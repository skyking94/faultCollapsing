module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,N425,N428,N429,N1fo0,N4fo0,N11fo0,N17fo0,N24fo0,N30fo0,N37fo0,N43fo0,N50fo0,N56fo0,N63fo0,N69fo0,N76fo0,N82fo0,N89fo0,N95fo0,N102fo0,N108fo0,N4fo1,N8fo0,N119fo0,N14fo0,N119fo1,N17fo1,N30fo1,N43fo1,N56fo1,N69fo1,N82fo1,N95fo1,N108fo1,N21fo0,N123fo0,N27fo0,N123fo1,N34fo0,N127fo0,N40fo0,N127fo1,N47fo0,N131fo0,N53fo0,N131fo1,N60fo0,N135fo0,N66fo0,N135fo1,N73fo0,N139fo0,N79fo0,N139fo1,N86fo0,N143fo0,N92fo0,N143fo1,N99fo0,N147fo0,N105fo0,N147fo1,N112fo0,N151fo0,N115fo0,N151fo1,N177fo0,N180fo0,N154fo0,N159fo0,N162fo0,N165fo0,N168fo0,N171fo0,N174fo0,N199fo0,N199fo1,N199fo2,N203fo0,N154fo1,N203fo1,N159fo1,N203fo2,N162fo1,N203fo3,N165fo1,N203fo4,N168fo1,N203fo5,N171fo1,N1fo1,N213fo0,N203fo6,N174fo1,N213fo1,N11fo1,N203fo7,N177fo1,N213fo2,N24fo1,N203fo8,N180fo1,N213fo3,N37fo1,N213fo4,N50fo1,N213fo5,N63fo1,N213fo6,N76fo1,N213fo7,N89fo1,N213fo8,N102fo1,N224fo0,N224fo1,N227fo0,N230fo0,N233fo0,N236fo0,N239fo0,N243fo0,N247fo0,N251fo0,N227fo1,N230fo1,N233fo1,N236fo1,N239fo1,N243fo1,N247fo1,N251fo1,N282fo0,N285fo0,N260fo0,N264fo0,N267fo0,N270fo0,N273fo0,N276fo0,N279fo0,N296fo0,N296fo1,N296fo2,N309fo0,N260fo1,N309fo1,N264fo1,N309fo2,N267fo1,N309fo3,N270fo1,N8fo1,N319fo0,N309fo4,N273fo1,N319fo1,N21fo1,N309fo5,N276fo1,N319fo2,N34fo1,N309fo6,N279fo1,N319fo3,N47fo1,N309fo7,N282fo1,N319fo4,N60fo1,N309fo8,N285fo1,N319fo5,N73fo1,N319fo6,N86fo1,N319fo7,N99fo1,N319fo8,N112fo1,N357fo0,N357fo1,N14fo1,N360fo0,N360fo1,N27fo1,N360fo2,N40fo1,N360fo3,N53fo1,N360fo4,N66fo1,N360fo5,N79fo1,N360fo6,N92fo1,N360fo7,N105fo1,N360fo8,N115fo1,N4fo2,N17fo2,N30fo2,N43fo2,N56fo2,N69fo2,N82fo2,N95fo2,N108fo2,N411fo0,N381fo0,N386fo0,N393fo0,N399fo0,N404fo0,N407fo0,N393fo1,N404fo1,N407fo1,N411fo1,N386fo1,N399fo1,N386fo2,N393fo2,N393fo3,N399fo2,N407fo2,N386fo3,N393fo4,N422fo0,N399fo3,N381fo1,N386fo4,N425fo0,N381fo2,N386fo5,N425fo1,N381fo3,N422fo1;
INVX1 uut0 (.Y(N118),.A(N1fo0));
INVX1 uut1 (.Y(N119),.A(N4fo0));
INVX1 uut2 (.Y(N122),.A(N11fo0));
INVX1 uut3 (.Y(N123),.A(N17fo0));
INVX1 uut4 (.Y(N126),.A(N24fo0));
INVX1 uut5 (.Y(N127),.A(N30fo0));
INVX1 uut6 (.Y(N130),.A(N37fo0));
INVX1 uut7 (.Y(N131),.A(N43fo0));
INVX1 uut8 (.Y(N134),.A(N50fo0));
INVX1 uut9 (.Y(N135),.A(N56fo0));
INVX1 uut10 (.Y(N138),.A(N63fo0));
INVX1 uut11 (.Y(N139),.A(N69fo0));
INVX1 uut12 (.Y(N142),.A(N76fo0));
INVX1 uut13 (.Y(N143),.A(N82fo0));
INVX1 uut14 (.Y(N146),.A(N89fo0));
INVX1 uut15 (.Y(N147),.A(N95fo0));
INVX1 uut16 (.Y(N150),.A(N102fo0));
INVX1 uut17 (.Y(N151),.A(N108fo0));
NAND2X1 uut18 (.Y(N154),.A(N118),.B(N4fo1));
NOR2X1 uut19 (.Y(N157),.A(N8fo0),.B(N119fo0));
NOR2X1 uut20 (.Y(N158),.A(N14fo0),.B(N119fo1));
NAND2X1 uut21 (.Y(N159),.A(N122),.B(N17fo1));
NAND2X1 uut22 (.Y(N162),.A(N126),.B(N30fo1));
NAND2X1 uut23 (.Y(N165),.A(N130),.B(N43fo1));
NAND2X1 uut24 (.Y(N168),.A(N134),.B(N56fo1));
NAND2X1 uut25 (.Y(N171),.A(N138),.B(N69fo1));
NAND2X1 uut26 (.Y(N174),.A(N142),.B(N82fo1));
NAND2X1 uut27 (.Y(N177),.A(N146),.B(N95fo1));
NAND2X1 uut28 (.Y(N180),.A(N150),.B(N108fo1));
NOR2X1 uut29 (.Y(N183),.A(N21fo0),.B(N123fo0));
NOR2X1 uut30 (.Y(N184),.A(N27fo0),.B(N123fo1));
NOR2X1 uut31 (.Y(N185),.A(N34fo0),.B(N127fo0));
NOR2X1 uut32 (.Y(N186),.A(N40fo0),.B(N127fo1));
NOR2X1 uut33 (.Y(N187),.A(N47fo0),.B(N131fo0));
NOR2X1 uut34 (.Y(N188),.A(N53fo0),.B(N131fo1));
NOR2X1 uut35 (.Y(N189),.A(N60fo0),.B(N135fo0));
NOR2X1 uut36 (.Y(N190),.A(N66fo0),.B(N135fo1));
NOR2X1 uut37 (.Y(N191),.A(N73fo0),.B(N139fo0));
NOR2X1 uut38 (.Y(N192),.A(N79fo0),.B(N139fo1));
NOR2X1 uut39 (.Y(N193),.A(N86fo0),.B(N143fo0));
NOR2X1 uut40 (.Y(N194),.A(N92fo0),.B(N143fo1));
NOR2X1 uut41 (.Y(N195),.A(N99fo0),.B(N147fo0));
NOR2X1 uut42 (.Y(N196),.A(N105fo0),.B(N147fo1));
NOR2X1 uut43 (.Y(N197),.A(N112fo0),.B(N151fo0));
NOR2X1 uut44 (.Y(N198),.A(N115fo0),.B(N151fo1));
AND2X1 uut45 (.Y(ttmp1),.A(N177fo0),.B(N180fo0));
AND2X1 uut46 (.Y(ttmp2),.A(N154fo0),.B(ttmp1));
AND2X1 uut47 (.Y(ttmp3),.A(N159fo0),.B(ttmp2));
AND2X1 uut48 (.Y(ttmp4),.A(N162fo0),.B(ttmp3));
AND2X1 uut49 (.Y(ttmp5),.A(N165fo0),.B(ttmp4));
AND2X1 uut50 (.Y(ttmp6),.A(N168fo0),.B(ttmp5));
AND2X1 uut51 (.Y(ttmp7),.A(N171fo0),.B(ttmp6));
AND2X1 uut52 (.Y(N199),.A(N174fo0),.B(ttmp7));
INVX1 uut53 (.Y(N203),.A(N199fo0));
INVX1 uut54 (.Y(N213),.A(N199fo1));
INVX1 uut55 (.Y(N223),.A(N199fo2));
XOR2X1 uut56 (.Y(N224),.A(N203fo0),.B(N154fo1));
XOR2X1 uut57 (.Y(N227),.A(N203fo1),.B(N159fo1));
XOR2X1 uut58 (.Y(N230),.A(N203fo2),.B(N162fo1));
XOR2X1 uut59 (.Y(N233),.A(N203fo3),.B(N165fo1));
XOR2X1 uut60 (.Y(N236),.A(N203fo4),.B(N168fo1));
XOR2X1 uut61 (.Y(N239),.A(N203fo5),.B(N171fo1));
NAND2X1 uut62 (.Y(N242),.A(N1fo1),.B(N213fo0));
XOR2X1 uut63 (.Y(N243),.A(N203fo6),.B(N174fo1));
NAND2X1 uut64 (.Y(N246),.A(N213fo1),.B(N11fo1));
XOR2X1 uut65 (.Y(N247),.A(N203fo7),.B(N177fo1));
NAND2X1 uut66 (.Y(N250),.A(N213fo2),.B(N24fo1));
XOR2X1 uut67 (.Y(N251),.A(N203fo8),.B(N180fo1));
NAND2X1 uut68 (.Y(N254),.A(N213fo3),.B(N37fo1));
NAND2X1 uut69 (.Y(N255),.A(N213fo4),.B(N50fo1));
NAND2X1 uut70 (.Y(N256),.A(N213fo5),.B(N63fo1));
NAND2X1 uut71 (.Y(N257),.A(N213fo6),.B(N76fo1));
NAND2X1 uut72 (.Y(N258),.A(N213fo7),.B(N89fo1));
NAND2X1 uut73 (.Y(N259),.A(N213fo8),.B(N102fo1));
NAND2X1 uut74 (.Y(N260),.A(N224fo0),.B(N157));
NAND2X1 uut75 (.Y(N263),.A(N224fo1),.B(N158));
NAND2X1 uut76 (.Y(N264),.A(N227fo0),.B(N183));
NAND2X1 uut77 (.Y(N267),.A(N230fo0),.B(N185));
NAND2X1 uut78 (.Y(N270),.A(N233fo0),.B(N187));
NAND2X1 uut79 (.Y(N273),.A(N236fo0),.B(N189));
NAND2X1 uut80 (.Y(N276),.A(N239fo0),.B(N191));
NAND2X1 uut81 (.Y(N279),.A(N243fo0),.B(N193));
NAND2X1 uut82 (.Y(N282),.A(N247fo0),.B(N195));
NAND2X1 uut83 (.Y(N285),.A(N251fo0),.B(N197));
NAND2X1 uut84 (.Y(N288),.A(N227fo1),.B(N184));
NAND2X1 uut85 (.Y(N289),.A(N230fo1),.B(N186));
NAND2X1 uut86 (.Y(N290),.A(N233fo1),.B(N188));
NAND2X1 uut87 (.Y(N291),.A(N236fo1),.B(N190));
NAND2X1 uut88 (.Y(N292),.A(N239fo1),.B(N192));
NAND2X1 uut89 (.Y(N293),.A(N243fo1),.B(N194));
NAND2X1 uut90 (.Y(N294),.A(N247fo1),.B(N196));
NAND2X1 uut91 (.Y(N295),.A(N251fo1),.B(N198));
AND2X1 uut92 (.Y(ttmp9),.A(N282fo0),.B(N285fo0));
AND2X1 uut93 (.Y(ttmp10),.A(N260fo0),.B(ttmp9));
AND2X1 uut94 (.Y(ttmp11),.A(N264fo0),.B(ttmp10));
AND2X1 uut95 (.Y(ttmp12),.A(N267fo0),.B(ttmp11));
AND2X1 uut96 (.Y(ttmp13),.A(N270fo0),.B(ttmp12));
AND2X1 uut97 (.Y(ttmp14),.A(N273fo0),.B(ttmp13));
AND2X1 uut98 (.Y(ttmp15),.A(N276fo0),.B(ttmp14));
AND2X1 uut99 (.Y(N296),.A(N279fo0),.B(ttmp15));
INVX1 uut100 (.Y(N300),.A(N263));
INVX1 uut101 (.Y(N301),.A(N288));
INVX1 uut102 (.Y(N302),.A(N289));
INVX1 uut103 (.Y(N303),.A(N290));
INVX1 uut104 (.Y(N304),.A(N291));
INVX1 uut105 (.Y(N305),.A(N292));
INVX1 uut106 (.Y(N306),.A(N293));
INVX1 uut107 (.Y(N307),.A(N294));
INVX1 uut108 (.Y(N308),.A(N295));
INVX1 uut109 (.Y(N309),.A(N296fo0));
INVX1 uut110 (.Y(N319),.A(N296fo1));
INVX1 uut111 (.Y(N329),.A(N296fo2));
XOR2X1 uut112 (.Y(N330),.A(N309fo0),.B(N260fo1));
XOR2X1 uut113 (.Y(N331),.A(N309fo1),.B(N264fo1));
XOR2X1 uut114 (.Y(N332),.A(N309fo2),.B(N267fo1));
XOR2X1 uut115 (.Y(N333),.A(N309fo3),.B(N270fo1));
NAND2X1 uut116 (.Y(N334),.A(N8fo1),.B(N319fo0));
XOR2X1 uut117 (.Y(N335),.A(N309fo4),.B(N273fo1));
NAND2X1 uut118 (.Y(N336),.A(N319fo1),.B(N21fo1));
XOR2X1 uut119 (.Y(N337),.A(N309fo5),.B(N276fo1));
NAND2X1 uut120 (.Y(N338),.A(N319fo2),.B(N34fo1));
XOR2X1 uut121 (.Y(N339),.A(N309fo6),.B(N279fo1));
NAND2X1 uut122 (.Y(N340),.A(N319fo3),.B(N47fo1));
XOR2X1 uut123 (.Y(N341),.A(N309fo7),.B(N282fo1));
NAND2X1 uut124 (.Y(N342),.A(N319fo4),.B(N60fo1));
XOR2X1 uut125 (.Y(N343),.A(N309fo8),.B(N285fo1));
NAND2X1 uut126 (.Y(N344),.A(N319fo5),.B(N73fo1));
NAND2X1 uut127 (.Y(N345),.A(N319fo6),.B(N86fo1));
NAND2X1 uut128 (.Y(N346),.A(N319fo7),.B(N99fo1));
NAND2X1 uut129 (.Y(N347),.A(N319fo8),.B(N112fo1));
NAND2X1 uut130 (.Y(N348),.A(N330),.B(N300));
NAND2X1 uut131 (.Y(N349),.A(N331),.B(N301));
NAND2X1 uut132 (.Y(N350),.A(N332),.B(N302));
NAND2X1 uut133 (.Y(N351),.A(N333),.B(N303));
NAND2X1 uut134 (.Y(N352),.A(N335),.B(N304));
NAND2X1 uut135 (.Y(N353),.A(N337),.B(N305));
NAND2X1 uut136 (.Y(N354),.A(N339),.B(N306));
NAND2X1 uut137 (.Y(N355),.A(N341),.B(N307));
NAND2X1 uut138 (.Y(N356),.A(N343),.B(N308));
AND2X1 uut139 (.Y(ttmp17),.A(N355),.B(N356));
AND2X1 uut140 (.Y(ttmp18),.A(N348),.B(ttmp17));
AND2X1 uut141 (.Y(ttmp19),.A(N349),.B(ttmp18));
AND2X1 uut142 (.Y(ttmp20),.A(N350),.B(ttmp19));
AND2X1 uut143 (.Y(ttmp21),.A(N351),.B(ttmp20));
AND2X1 uut144 (.Y(ttmp22),.A(N352),.B(ttmp21));
AND2X1 uut145 (.Y(ttmp23),.A(N353),.B(ttmp22));
AND2X1 uut146 (.Y(N357),.A(N354),.B(ttmp23));
INVX1 uut147 (.Y(N360),.A(N357fo0));
INVX1 uut148 (.Y(N370),.A(N357fo1));
NAND2X1 uut149 (.Y(N371),.A(N14fo1),.B(N360fo0));
NAND2X1 uut150 (.Y(N372),.A(N360fo1),.B(N27fo1));
NAND2X1 uut151 (.Y(N373),.A(N360fo2),.B(N40fo1));
NAND2X1 uut152 (.Y(N374),.A(N360fo3),.B(N53fo1));
NAND2X1 uut153 (.Y(N375),.A(N360fo4),.B(N66fo1));
NAND2X1 uut154 (.Y(N376),.A(N360fo5),.B(N79fo1));
NAND2X1 uut155 (.Y(N377),.A(N360fo6),.B(N92fo1));
NAND2X1 uut156 (.Y(N378),.A(N360fo7),.B(N105fo1));
NAND2X1 uut157 (.Y(N379),.A(N360fo8),.B(N115fo1));
AND2X1 uut158 (.Y(ttmp25),.A(N334),.B(N371));
AND2X1 uut159 (.Y(ttmp26),.A(N4fo2),.B(ttmp25));
NAND2X1 uut160 (.Y(N380),.A(N242),.B(ttmp26));
AND2X1 uut161 (.Y(ttmp28),.A(N372),.B(N17fo2));
AND2X1 uut162 (.Y(ttmp29),.A(N246),.B(ttmp28));
NAND2X1 uut163 (.Y(N381),.A(N336),.B(ttmp29));
AND2X1 uut164 (.Y(ttmp31),.A(N373),.B(N30fo2));
AND2X1 uut165 (.Y(ttmp32),.A(N250),.B(ttmp31));
NAND2X1 uut166 (.Y(N386),.A(N338),.B(ttmp32));
AND2X1 uut167 (.Y(ttmp34),.A(N374),.B(N43fo2));
AND2X1 uut168 (.Y(ttmp35),.A(N254),.B(ttmp34));
NAND2X1 uut169 (.Y(N393),.A(N340),.B(ttmp35));
AND2X1 uut170 (.Y(ttmp37),.A(N375),.B(N56fo2));
AND2X1 uut171 (.Y(ttmp38),.A(N255),.B(ttmp37));
NAND2X1 uut172 (.Y(N399),.A(N342),.B(ttmp38));
AND2X1 uut173 (.Y(ttmp40),.A(N376),.B(N69fo2));
AND2X1 uut174 (.Y(ttmp41),.A(N256),.B(ttmp40));
NAND2X1 uut175 (.Y(N404),.A(N344),.B(ttmp41));
AND2X1 uut176 (.Y(ttmp43),.A(N377),.B(N82fo2));
AND2X1 uut177 (.Y(ttmp44),.A(N257),.B(ttmp43));
NAND2X1 uut178 (.Y(N407),.A(N345),.B(ttmp44));
AND2X1 uut179 (.Y(ttmp46),.A(N378),.B(N95fo2));
AND2X1 uut180 (.Y(ttmp47),.A(N258),.B(ttmp46));
NAND2X1 uut181 (.Y(N411),.A(N346),.B(ttmp47));
AND2X1 uut182 (.Y(ttmp49),.A(N379),.B(N108fo2));
AND2X1 uut183 (.Y(ttmp50),.A(N259),.B(ttmp49));
NAND2X1 uut184 (.Y(N414),.A(N347),.B(ttmp50));
INVX1 uut185 (.Y(N415),.A(N380));
AND2X1 uut186 (.Y(ttmp52),.A(N411fo0),.B(N414));
AND2X1 uut187 (.Y(ttmp53),.A(N381fo0),.B(ttmp52));
AND2X1 uut188 (.Y(ttmp54),.A(N386fo0),.B(ttmp53));
AND2X1 uut189 (.Y(ttmp55),.A(N393fo0),.B(ttmp54));
AND2X1 uut190 (.Y(ttmp56),.A(N399fo0),.B(ttmp55));
AND2X1 uut191 (.Y(ttmp57),.A(N404fo0),.B(ttmp56));
AND2X1 uut192 (.Y(N416),.A(N407fo0),.B(ttmp57));
INVX1 uut193 (.Y(N417),.A(N393fo1));
INVX1 uut194 (.Y(N418),.A(N404fo1));
INVX1 uut195 (.Y(N419),.A(N407fo1));
INVX1 uut196 (.Y(N420),.A(N411fo1));
NOR2X1 uut197 (.Y(N421),.A(N415),.B(N416));
NAND2X1 uut198 (.Y(N422),.A(N386fo1),.B(N417));
AND2X1 uut199 (.Y(ttmp59),.A(N418),.B(N399fo1));
AND2X1 uut200 (.Y(ttmp60),.A(N386fo2),.B(ttmp59));
NAND2X1 uut201 (.Y(N425),.A(N393fo2),.B(ttmp60));
AND2X1 uut202 (.Y(ttmp62),.A(N393fo3),.B(N419));
NAND2X1 uut203 (.Y(N428),.A(N399fo2),.B(ttmp62));
AND2X1 uut204 (.Y(ttmp64),.A(N407fo2),.B(N420));
AND2X1 uut205 (.Y(ttmp65),.A(N386fo3),.B(ttmp64));
NAND2X1 uut206 (.Y(N429),.A(N393fo4),.B(ttmp65));
AND2X1 uut207 (.Y(ttmp67),.A(N422fo0),.B(N399fo3));
AND2X1 uut208 (.Y(ttmp68),.A(N381fo1),.B(ttmp67));
NAND2X1 uut209 (.Y(N430),.A(N386fo4),.B(ttmp68));
AND2X1 uut210 (.Y(ttmp70),.A(N425fo0),.B(N428));
AND2X1 uut211 (.Y(ttmp71),.A(N381fo2),.B(ttmp70));
NAND2X1 uut212 (.Y(N431),.A(N386fo5),.B(ttmp71));
AND2X1 uut213 (.Y(ttmp73),.A(N425fo1),.B(N429));
AND2X1 uut214 (.Y(ttmp74),.A(N381fo3),.B(ttmp73));
NAND2X1 uut215 (.Y(N432),.A(N422fo1),.B(ttmp74));
fanout2 uut_fo0 (.A(N1),.Y1(N1fo0),.Y2(N1fo1));
fanout3 uut_fo1 (.A(N4),.Y1(N4fo0),.Y2(N4fo1),.Y3(N4fo2));
fanout2 uut_fo2 (.A(N8),.Y1(N8fo0),.Y2(N8fo1));
fanout2 uut_fo3 (.A(N11),.Y1(N11fo0),.Y2(N11fo1));
fanout2 uut_fo4 (.A(N14),.Y1(N14fo0),.Y2(N14fo1));
fanout3 uut_fo5 (.A(N17),.Y1(N17fo0),.Y2(N17fo1),.Y3(N17fo2));
fanout2 uut_fo6 (.A(N21),.Y1(N21fo0),.Y2(N21fo1));
fanout2 uut_fo7 (.A(N24),.Y1(N24fo0),.Y2(N24fo1));
fanout2 uut_fo8 (.A(N27),.Y1(N27fo0),.Y2(N27fo1));
fanout3 uut_fo9 (.A(N30),.Y1(N30fo0),.Y2(N30fo1),.Y3(N30fo2));
fanout2 uut_fo10 (.A(N34),.Y1(N34fo0),.Y2(N34fo1));
fanout2 uut_fo11 (.A(N37),.Y1(N37fo0),.Y2(N37fo1));
fanout2 uut_fo12 (.A(N40),.Y1(N40fo0),.Y2(N40fo1));
fanout3 uut_fo13 (.A(N43),.Y1(N43fo0),.Y2(N43fo1),.Y3(N43fo2));
fanout2 uut_fo14 (.A(N47),.Y1(N47fo0),.Y2(N47fo1));
fanout2 uut_fo15 (.A(N50),.Y1(N50fo0),.Y2(N50fo1));
fanout2 uut_fo16 (.A(N53),.Y1(N53fo0),.Y2(N53fo1));
fanout3 uut_fo17 (.A(N56),.Y1(N56fo0),.Y2(N56fo1),.Y3(N56fo2));
fanout2 uut_fo18 (.A(N60),.Y1(N60fo0),.Y2(N60fo1));
fanout2 uut_fo19 (.A(N63),.Y1(N63fo0),.Y2(N63fo1));
fanout2 uut_fo20 (.A(N66),.Y1(N66fo0),.Y2(N66fo1));
fanout3 uut_fo21 (.A(N69),.Y1(N69fo0),.Y2(N69fo1),.Y3(N69fo2));
fanout2 uut_fo22 (.A(N73),.Y1(N73fo0),.Y2(N73fo1));
fanout2 uut_fo23 (.A(N76),.Y1(N76fo0),.Y2(N76fo1));
fanout2 uut_fo24 (.A(N79),.Y1(N79fo0),.Y2(N79fo1));
fanout3 uut_fo25 (.A(N82),.Y1(N82fo0),.Y2(N82fo1),.Y3(N82fo2));
fanout2 uut_fo26 (.A(N86),.Y1(N86fo0),.Y2(N86fo1));
fanout2 uut_fo27 (.A(N89),.Y1(N89fo0),.Y2(N89fo1));
fanout2 uut_fo28 (.A(N92),.Y1(N92fo0),.Y2(N92fo1));
fanout3 uut_fo29 (.A(N95),.Y1(N95fo0),.Y2(N95fo1),.Y3(N95fo2));
fanout2 uut_fo30 (.A(N99),.Y1(N99fo0),.Y2(N99fo1));
fanout2 uut_fo31 (.A(N102),.Y1(N102fo0),.Y2(N102fo1));
fanout2 uut_fo32 (.A(N105),.Y1(N105fo0),.Y2(N105fo1));
fanout3 uut_fo33 (.A(N108),.Y1(N108fo0),.Y2(N108fo1),.Y3(N108fo2));
fanout2 uut_fo34 (.A(N112),.Y1(N112fo0),.Y2(N112fo1));
fanout2 uut_fo35 (.A(N115),.Y1(N115fo0),.Y2(N115fo1));
fanout2 uut_fo_w0 (.A(N276),.Y1(N276fo0),.Y2(N276fo1));
fanout2 uut_fo_w1 (.A(N135),.Y1(N135fo0),.Y2(N135fo1));
fanout2 uut_fo_w15 (.A(N177),.Y1(N177fo0),.Y2(N177fo1));
fanout9 uut_fo_w20 (.A(N360),.Y1(N360fo0),.Y2(N360fo1),.Y3(N360fo2),.Y4(N360fo3),.Y5(N360fo4),.Y6(N360fo5),.Y7(N360fo6),.Y8(N360fo7),.Y9(N360fo8));
fanout2 uut_fo_w25 (.A(N279),.Y1(N279fo0),.Y2(N279fo1));
fanout2 uut_fo_w27 (.A(N174),.Y1(N174fo0),.Y2(N174fo1));
fanout9 uut_fo_w29 (.A(N203),.Y1(N203fo0),.Y2(N203fo1),.Y3(N203fo2),.Y4(N203fo3),.Y5(N203fo4),.Y6(N203fo5),.Y7(N203fo6),.Y8(N203fo7),.Y9(N203fo8));
fanout2 uut_fo_w31 (.A(N171),.Y1(N171fo0),.Y2(N171fo1));
fanout2 uut_fo_w44 (.A(N131),.Y1(N131fo0),.Y2(N131fo1));
fanout2 uut_fo_w45 (.A(N154),.Y1(N154fo0),.Y2(N154fo1));
fanout2 uut_fo_w46 (.A(N357),.Y1(N357fo0),.Y2(N357fo1));
fanout2 uut_fo_w48 (.A(N168),.Y1(N168fo0),.Y2(N168fo1));
fanout2 uut_fo_w51 (.A(N267),.Y1(N267fo0),.Y2(N267fo1));
fanout2 uut_fo_w57 (.A(N127),.Y1(N127fo0),.Y2(N127fo1));
fanout2 uut_fo_w59 (.A(N251),.Y1(N251fo0),.Y2(N251fo1));
fanout2 uut_fo_w63 (.A(N282),.Y1(N282fo0),.Y2(N282fo1));
fanout2 uut_fo_w64 (.A(N243),.Y1(N243fo0),.Y2(N243fo1));
fanout2 uut_fo_w67 (.A(N180),.Y1(N180fo0),.Y2(N180fo1));
fanout3 uut_fo_w73 (.A(N199),.Y1(N199fo0),.Y2(N199fo1),.Y3(N199fo2));
fanout2 uut_fo_w74 (.A(N422),.Y1(N422fo0),.Y2(N422fo1));
fanout2 uut_fo_w76 (.A(N411),.Y1(N411fo0),.Y2(N411fo1));
fanout2 uut_fo_w81 (.A(N224),.Y1(N224fo0),.Y2(N224fo1));
fanout2 uut_fo_w82 (.A(N285),.Y1(N285fo0),.Y2(N285fo1));
fanout2 uut_fo_w84 (.A(N139),.Y1(N139fo0),.Y2(N139fo1));
fanout2 uut_fo_w88 (.A(N159),.Y1(N159fo0),.Y2(N159fo1));
fanout2 uut_fo_w98 (.A(N162),.Y1(N162fo0),.Y2(N162fo1));
fanout2 uut_fo_w102 (.A(N227),.Y1(N227fo0),.Y2(N227fo1));
fanout2 uut_fo_w105 (.A(N143),.Y1(N143fo0),.Y2(N143fo1));
fanout9 uut_fo_w106 (.A(N309),.Y1(N309fo0),.Y2(N309fo1),.Y3(N309fo2),.Y4(N309fo3),.Y5(N309fo4),.Y6(N309fo5),.Y7(N309fo6),.Y8(N309fo7),.Y9(N309fo8));
fanout2 uut_fo_w109 (.A(N270),.Y1(N270fo0),.Y2(N270fo1));
fanout2 uut_fo_w110 (.A(N230),.Y1(N230fo0),.Y2(N230fo1));
fanout2 uut_fo_w121 (.A(N425),.Y1(N425fo0),.Y2(N425fo1));
fanout4 uut_fo_w130 (.A(N381),.Y1(N381fo0),.Y2(N381fo1),.Y3(N381fo2),.Y4(N381fo3));
fanout3 uut_fo_w132 (.A(N296),.Y1(N296fo0),.Y2(N296fo1),.Y3(N296fo2));
fanout2 uut_fo_w137 (.A(N165),.Y1(N165fo0),.Y2(N165fo1));
fanout9 uut_fo_w139 (.A(N213),.Y1(N213fo0),.Y2(N213fo1),.Y3(N213fo2),.Y4(N213fo3),.Y5(N213fo4),.Y6(N213fo5),.Y7(N213fo6),.Y8(N213fo7),.Y9(N213fo8));
fanout2 uut_fo_w144 (.A(N273),.Y1(N273fo0),.Y2(N273fo1));
fanout2 uut_fo_w148 (.A(N239),.Y1(N239fo0),.Y2(N239fo1));
fanout5 uut_fo_w149 (.A(N393),.Y1(N393fo0),.Y2(N393fo1),.Y3(N393fo2),.Y4(N393fo3),.Y5(N393fo4));
fanout2 uut_fo_w152 (.A(N404),.Y1(N404fo0),.Y2(N404fo1));
fanout2 uut_fo_w159 (.A(N260),.Y1(N260fo0),.Y2(N260fo1));
fanout2 uut_fo_w168 (.A(N147),.Y1(N147fo0),.Y2(N147fo1));
fanout2 uut_fo_w169 (.A(N233),.Y1(N233fo0),.Y2(N233fo1));
fanout6 uut_fo_w170 (.A(N386),.Y1(N386fo0),.Y2(N386fo1),.Y3(N386fo2),.Y4(N386fo3),.Y5(N386fo4),.Y6(N386fo5));
fanout2 uut_fo_w171 (.A(N247),.Y1(N247fo0),.Y2(N247fo1));
fanout9 uut_fo_w177 (.A(N319),.Y1(N319fo0),.Y2(N319fo1),.Y3(N319fo2),.Y4(N319fo3),.Y5(N319fo4),.Y6(N319fo5),.Y7(N319fo6),.Y8(N319fo7),.Y9(N319fo8));
fanout2 uut_fo_w180 (.A(N236),.Y1(N236fo0),.Y2(N236fo1));
fanout2 uut_fo_w184 (.A(N123),.Y1(N123fo0),.Y2(N123fo1));
fanout2 uut_fo_w186 (.A(N264),.Y1(N264fo0),.Y2(N264fo1));
fanout2 uut_fo_w188 (.A(N151),.Y1(N151fo0),.Y2(N151fo1));
fanout3 uut_fo_w200 (.A(N407),.Y1(N407fo0),.Y2(N407fo1),.Y3(N407fo2));
fanout4 uut_fo_w202 (.A(N399),.Y1(N399fo0),.Y2(N399fo1),.Y3(N399fo2),.Y4(N399fo3));
fanout2 uut_fo_w207 (.A(N119),.Y1(N119fo0),.Y2(N119fo1));
endmodule