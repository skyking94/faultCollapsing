module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,N870,N871,N872,N873,N875,N876,N877,N13fo0,N17fo0,N1fo0,N8fo0,N13fo1,N17fo1,N1fo1,N26fo0,N36fo0,N42fo0,N29fo0,N26fo1,N51fo0,N1fo2,N51fo1,N17fo2,N1fo3,N8fo1,N13fo2,N55fo0,N1fo4,N8fo2,N68fo0,N59fo0,N42fo1,N29fo1,N68fo1,N68fo2,N59fo1,N75fo0,N80fo0,N29fo2,N75fo1,N42fo2,N29fo3,N36fo1,N80fo1,N29fo4,N36fo2,N42fo3,N29fo5,N75fo2,N80fo2,N59fo2,N75fo3,N42fo4,N59fo3,N36fo3,N80fo3,N59fo4,N36fo4,N42fo5,N59fo5,N91fo0,N96fo0,N91fo1,N96fo1,N101fo0,N106fo0,N101fo1,N106fo1,N111fo0,N116fo0,N111fo1,N116fo1,N121fo0,N126fo0,N121fo1,N126fo1,N8fo3,N138fo0,N51fo2,N138fo1,N17fo3,N138fo2,N138fo3,N59fo6,N156fo0,N17fo4,N42fo6,N17fo5,N42fo7,N159fo0,N165fo0,N159fo1,N165fo1,N171fo0,N177fo0,N171fo1,N177fo1,N183fo0,N189fo0,N183fo1,N189fo1,N195fo0,N201fo0,N195fo1,N201fo1,N210fo0,N91fo2,N210fo1,N96fo2,N210fo2,N101fo2,N210fo3,N106fo2,N210fo4,N111fo2,N255fo0,N210fo5,N116fo2,N255fo1,N210fo6,N121fo2,N255fo2,N273fo0,N270fo0,N273fo1,N276fo0,N276fo1,N280fo0,N280fo1,N280fo2,N298fo0,N298fo1,N310fo0,N270fo1,N357fo0,N360fo0,N357fo1,N360fo1,N363fo0,N366fo0,N363fo1,N366fo1,N376fo0,N379fo0,N376fo1,N379fo1,N382fo0,N385fo0,N382fo1,N385fo1,N210fo7,N369fo0,N393fo0,N55fo1,N319fo0,N17fo6,N287fo0,N393fo1,N287fo1,N55fo2,N393fo2,N156fo1,N393fo3,N59fo7,N319fo1,N17fo7,N393fo4,N143fo0,N427fo0,N310fo1,N432fo0,N146fo0,N427fo1,N310fo2,N432fo1,N149fo0,N427fo2,N310fo3,N432fo2,N153fo0,N427fo3,N310fo4,N432fo3,N1fo5,N369fo1,N437fo0,N369fo2,N437fo1,N369fo3,N437fo2,N369fo4,N437fo3,N130fo0,N460fo0,N130fo1,N460fo1,N463fo0,N135fo0,N463fo1,N135fo1,N91fo3,N466fo0,N96fo3,N466fo1,N101fo3,N466fo2,N106fo3,N466fo3,N143fo1,N483fo0,N111fo3,N466fo4,N146fo1,N483fo1,N116fo3,N466fo5,N149fo1,N483fo2,N121fo3,N466fo6,N153fo1,N483fo3,N126fo2,N466fo7,N130fo2,N492fo0,N130fo3,N492fo1,N495fo0,N207fo0,N495fo1,N207fo1,N451fo0,N159fo2,N451fo1,N165fo2,N451fo2,N171fo2,N451fo3,N177fo2,N451fo4,N183fo2,N451fo5,N189fo2,N451fo6,N195fo2,N451fo7,N201fo2,N530fo0,N533fo0,N530fo1,N533fo1,N544fo0,N547fo0,N544fo1,N547fo1,N553fo0,N159fo3,N553fo1,N159fo4,N246fo0,N553fo2,N557fo0,N165fo3,N557fo1,N165fo4,N246fo1,N557fo2,N561fo0,N171fo3,N561fo1,N171fo4,N246fo2,N561fo2,N565fo0,N177fo3,N565fo1,N177fo4,N246fo3,N565fo2,N569fo0,N183fo3,N569fo1,N183fo4,N246fo4,N569fo2,N573fo0,N189fo3,N573fo1,N189fo4,N246fo5,N573fo2,N577fo0,N195fo3,N577fo1,N195fo4,N246fo6,N577fo2,N581fo0,N201fo3,N581fo1,N201fo4,N246fo7,N581fo2,N590fo0,N593fo0,N590fo1,N597fo0,N600fo0,N597fo1,N606fo0,N609fo0,N606fo1,N616fo0,N619fo0,N616fo1,N625fo0,N628fo0,N625fo1,N632fo0,N635fo0,N632fo1,N641fo0,N644fo0,N641fo1,N651fo0,N654fo0,N651fo1,N654fo1,N261fo0,N654fo2,N261fo1,N644fo1,N654fo3,N261fo2,N635fo1,N644fo2,N662fo0,N228fo0,N665fo0,N237fo0,N662fo1,N670fo0,N228fo1,N673fo0,N237fo1,N670fo1,N678fo0,N228fo2,N682fo0,N237fo2,N678fo1,N687fo0,N228fo3,N692fo0,N237fo3,N687fo1,N697fo0,N228fo4,N700fo0,N237fo4,N697fo1,N705fo0,N228fo5,N708fo0,N237fo5,N705fo1,N713fo0,N228fo6,N717fo0,N237fo6,N713fo1,N722fo0,N727fo0,N261fo3,N727fo1,N261fo4,N228fo7,N727fo2,N237fo7,N722fo1,N644fo3,N722fo2,N635fo2,N713fo2,N644fo4,N722fo3,N635fo3,N609fo1,N687fo2,N600fo1,N678fo2,N609fo2,N687fo3,N600fo2,N700fo1,N773fo0,N700fo2,N773fo1,N708fo1,N778fo0,N708fo2,N778fo1,N717fo1,N782fo0,N717fo2,N782fo1,N219fo0,N628fo1,N773fo2,N692fo1,N796fo0,N692fo2,N796fo1,N219fo1,N219fo2,N219fo3,N619fo1,N796fo2,N619fo2,N796fo3,N609fo3,N619fo3,N796fo4,N600fo3,N609fo4,N665fo1,N815fo0,N665fo2,N815fo1,N673fo1,N819fo0,N673fo2,N819fo1,N682fo1,N822fo0,N682fo2,N822fo1,N219fo4,N815fo2,N593fo1,N219fo5,N219fo6,N219fo7;
AND2X1 uut0 (.Y(ttmp1),.A(N13fo0),.B(N17fo0));
AND2X1 uut1 (.Y(ttmp2),.A(N1fo0),.B(ttmp1));
NAND2X1 uut2 (.Y(N269),.A(N8fo0),.B(ttmp2));
AND2X1 uut3 (.Y(ttmp4),.A(N13fo1),.B(N17fo1));
AND2X1 uut4 (.Y(ttmp5),.A(N1fo1),.B(ttmp4));
NAND2X1 uut5 (.Y(N270),.A(N26fo0),.B(ttmp5));
AND2X1 uut6 (.Y(ttmp7),.A(N36fo0),.B(N42fo0));
AND2X1 uut7 (.Y(N273),.A(N29fo0),.B(ttmp7));
AND2X1 uut8 (.Y(ttmp9),.A(N26fo1),.B(N51fo0));
AND2X1 uut9 (.Y(N276),.A(N1fo2),.B(ttmp9));
AND2X1 uut10 (.Y(ttmp11),.A(N51fo1),.B(N17fo2));
AND2X1 uut11 (.Y(ttmp12),.A(N1fo3),.B(ttmp11));
NAND2X1 uut12 (.Y(N279),.A(N8fo1),.B(ttmp12));
AND2X1 uut13 (.Y(ttmp14),.A(N13fo2),.B(N55fo0));
AND2X1 uut14 (.Y(ttmp15),.A(N1fo4),.B(ttmp14));
NAND2X1 uut15 (.Y(N280),.A(N8fo2),.B(ttmp15));
AND2X1 uut16 (.Y(ttmp17),.A(N68fo0),.B(N72));
AND2X1 uut17 (.Y(ttmp18),.A(N59fo0),.B(ttmp17));
NAND2X1 uut18 (.Y(N284),.A(N42fo1),.B(ttmp18));
NAND2X1 uut19 (.Y(N285),.A(N29fo1),.B(N68fo1));
AND2X1 uut20 (.Y(ttmp20),.A(N68fo2),.B(N74));
NAND2X1 uut21 (.Y(N286),.A(N59fo1),.B(ttmp20));
AND2X1 uut22 (.Y(ttmp22),.A(N75fo0),.B(N80fo0));
AND2X1 uut23 (.Y(N287),.A(N29fo2),.B(ttmp22));
AND2X1 uut24 (.Y(ttmp24),.A(N75fo1),.B(N42fo2));
AND2X1 uut25 (.Y(N290),.A(N29fo3),.B(ttmp24));
AND2X1 uut26 (.Y(ttmp26),.A(N36fo1),.B(N80fo1));
AND2X1 uut27 (.Y(N291),.A(N29fo4),.B(ttmp26));
AND2X1 uut28 (.Y(ttmp28),.A(N36fo2),.B(N42fo3));
AND2X1 uut29 (.Y(N292),.A(N29fo5),.B(ttmp28));
AND2X1 uut30 (.Y(ttmp30),.A(N75fo2),.B(N80fo2));
AND2X1 uut31 (.Y(N293),.A(N59fo2),.B(ttmp30));
AND2X1 uut32 (.Y(ttmp32),.A(N75fo3),.B(N42fo4));
AND2X1 uut33 (.Y(N294),.A(N59fo3),.B(ttmp32));
AND2X1 uut34 (.Y(ttmp34),.A(N36fo3),.B(N80fo3));
AND2X1 uut35 (.Y(N295),.A(N59fo4),.B(ttmp34));
AND2X1 uut36 (.Y(ttmp36),.A(N36fo4),.B(N42fo5));
AND2X1 uut37 (.Y(N296),.A(N59fo5),.B(ttmp36));
AND2X1 uut38 (.Y(N297),.A(N85),.B(N86));
OR2X1 uut39 (.Y(N298),.A(N87),.B(N88));
NAND2X1 uut40 (.Y(N301),.A(N91fo0),.B(N96fo0));
OR2X1 uut41 (.Y(N302),.A(N91fo1),.B(N96fo1));
NAND2X1 uut42 (.Y(N303),.A(N101fo0),.B(N106fo0));
OR2X1 uut43 (.Y(N304),.A(N101fo1),.B(N106fo1));
NAND2X1 uut44 (.Y(N305),.A(N111fo0),.B(N116fo0));
OR2X1 uut45 (.Y(N306),.A(N111fo1),.B(N116fo1));
NAND2X1 uut46 (.Y(N307),.A(N121fo0),.B(N126fo0));
OR2X1 uut47 (.Y(N308),.A(N121fo1),.B(N126fo1));
AND2X1 uut48 (.Y(N309),.A(N8fo3),.B(N138fo0));
INVX1 uut49 (.Y(N310),.A(N268));
AND2X1 uut50 (.Y(N316),.A(N51fo2),.B(N138fo1));
AND2X1 uut51 (.Y(N317),.A(N17fo3),.B(N138fo2));
AND2X1 uut52 (.Y(N318),.A(N152),.B(N138fo3));
NAND2X1 uut53 (.Y(N319),.A(N59fo6),.B(N156fo0));
NOR2X1 uut54 (.Y(N322),.A(N17fo4),.B(N42fo6));
AND2X1 uut55 (.Y(N323),.A(N17fo5),.B(N42fo7));
NAND2X1 uut56 (.Y(N324),.A(N159fo0),.B(N165fo0));
OR2X1 uut57 (.Y(N325),.A(N159fo1),.B(N165fo1));
NAND2X1 uut58 (.Y(N326),.A(N171fo0),.B(N177fo0));
OR2X1 uut59 (.Y(N327),.A(N171fo1),.B(N177fo1));
NAND2X1 uut60 (.Y(N328),.A(N183fo0),.B(N189fo0));
OR2X1 uut61 (.Y(N329),.A(N183fo1),.B(N189fo1));
NAND2X1 uut62 (.Y(N330),.A(N195fo0),.B(N201fo0));
OR2X1 uut63 (.Y(N331),.A(N195fo1),.B(N201fo1));
AND2X1 uut64 (.Y(N332),.A(N210fo0),.B(N91fo2));
AND2X1 uut65 (.Y(N333),.A(N210fo1),.B(N96fo2));
AND2X1 uut66 (.Y(N334),.A(N210fo2),.B(N101fo2));
AND2X1 uut67 (.Y(N335),.A(N210fo3),.B(N106fo2));
AND2X1 uut68 (.Y(N336),.A(N210fo4),.B(N111fo2));
AND2X1 uut69 (.Y(N337),.A(N255fo0),.B(N259));
AND2X1 uut70 (.Y(N338),.A(N210fo5),.B(N116fo2));
AND2X1 uut71 (.Y(N339),.A(N255fo1),.B(N260));
AND2X1 uut72 (.Y(N340),.A(N210fo6),.B(N121fo2));
AND2X1 uut73 (.Y(N341),.A(N255fo2),.B(N267));
INVX1 uut74 (.Y(N342),.A(N269));
INVX1 uut75 (.Y(N343),.A(N273fo0));
OR2X1 uut76 (.Y(N344),.A(N270fo0),.B(N273fo1));
INVX1 uut77 (.Y(N345),.A(N276fo0));
INVX1 uut78 (.Y(N346),.A(N276fo1));
INVX1 uut79 (.Y(N347),.A(N279));
NOR2X1 uut80 (.Y(N348),.A(N280fo0),.B(N284));
OR2X1 uut81 (.Y(N349),.A(N280fo1),.B(N285));
OR2X1 uut82 (.Y(N350),.A(N280fo2),.B(N286));
INVX1 uut83 (.Y(N351),.A(N293));
INVX1 uut84 (.Y(N352),.A(N294));
INVX1 uut85 (.Y(N353),.A(N295));
INVX1 uut86 (.Y(N354),.A(N296));
NAND2X1 uut87 (.Y(N355),.A(N89),.B(N298fo0));
AND2X1 uut88 (.Y(N356),.A(N90),.B(N298fo1));
NAND2X1 uut89 (.Y(N357),.A(N301),.B(N302));
NAND2X1 uut90 (.Y(N360),.A(N303),.B(N304));
NAND2X1 uut91 (.Y(N363),.A(N305),.B(N306));
NAND2X1 uut92 (.Y(N366),.A(N307),.B(N308));
INVX1 uut93 (.Y(N369),.A(N310fo0));
NOR2X1 uut94 (.Y(N375),.A(N322),.B(N323));
NAND2X1 uut95 (.Y(N376),.A(N324),.B(N325));
NAND2X1 uut96 (.Y(N379),.A(N326),.B(N327));
NAND2X1 uut97 (.Y(N382),.A(N328),.B(N329));
NAND2X1 uut98 (.Y(N385),.A(N330),.B(N331));
BUFX1 uut99 (.Y(N388),.A(N290));
BUFX1 uut100 (.Y(N389),.A(N291));
BUFX1 uut101 (.Y(N390),.A(N292));
BUFX1 uut102 (.Y(N391),.A(N297));
OR2X1 uut103 (.Y(N392),.A(N270fo1),.B(N343));
INVX1 uut104 (.Y(N393),.A(N345));
INVX1 uut105 (.Y(N399),.A(N346));
AND2X1 uut106 (.Y(N400),.A(N348),.B(N73));
INVX1 uut107 (.Y(N401),.A(N349));
INVX1 uut108 (.Y(N402),.A(N350));
INVX1 uut109 (.Y(N403),.A(N355));
INVX1 uut110 (.Y(N404),.A(N357fo0));
INVX1 uut111 (.Y(N405),.A(N360fo0));
AND2X1 uut112 (.Y(N406),.A(N357fo1),.B(N360fo1));
INVX1 uut113 (.Y(N407),.A(N363fo0));
INVX1 uut114 (.Y(N408),.A(N366fo0));
AND2X1 uut115 (.Y(N409),.A(N363fo1),.B(N366fo1));
NAND2X1 uut116 (.Y(N410),.A(N347),.B(N352));
INVX1 uut117 (.Y(N411),.A(N376fo0));
INVX1 uut118 (.Y(N412),.A(N379fo0));
AND2X1 uut119 (.Y(N413),.A(N376fo1),.B(N379fo1));
INVX1 uut120 (.Y(N414),.A(N382fo0));
INVX1 uut121 (.Y(N415),.A(N385fo0));
AND2X1 uut122 (.Y(N416),.A(N382fo1),.B(N385fo1));
AND2X1 uut123 (.Y(N417),.A(N210fo7),.B(N369fo0));
BUFX1 uut124 (.Y(N418),.A(N342));
BUFX1 uut125 (.Y(N419),.A(N344));
BUFX1 uut126 (.Y(N420),.A(N351));
BUFX1 uut127 (.Y(N421),.A(N353));
BUFX1 uut128 (.Y(N422),.A(N354));
BUFX1 uut129 (.Y(N423),.A(N356));
INVX1 uut130 (.Y(N424),.A(N400));
AND2X1 uut131 (.Y(N425),.A(N404),.B(N405));
AND2X1 uut132 (.Y(N426),.A(N407),.B(N408));
AND2X1 uut133 (.Y(ttmp38),.A(N393fo0),.B(N55fo1));
AND2X1 uut134 (.Y(N427),.A(N319fo0),.B(ttmp38));
AND2X1 uut135 (.Y(ttmp40),.A(N17fo6),.B(N287fo0));
AND2X1 uut136 (.Y(N432),.A(N393fo1),.B(ttmp40));
AND2X1 uut137 (.Y(ttmp42),.A(N287fo1),.B(N55fo2));
NAND2X1 uut138 (.Y(N437),.A(N393fo2),.B(ttmp42));
AND2X1 uut139 (.Y(ttmp44),.A(N156fo1),.B(N393fo3));
AND2X1 uut140 (.Y(ttmp45),.A(N375),.B(ttmp44));
NAND2X1 uut141 (.Y(N442),.A(N59fo7),.B(ttmp45));
AND2X1 uut142 (.Y(ttmp47),.A(N319fo1),.B(N17fo7));
NAND2X1 uut143 (.Y(N443),.A(N393fo4),.B(ttmp47));
AND2X1 uut144 (.Y(N444),.A(N411),.B(N412));
AND2X1 uut145 (.Y(N445),.A(N414),.B(N415));
BUFX1 uut146 (.Y(N446),.A(N392));
BUFX1 uut147 (.Y(N447),.A(N399));
BUFX1 uut148 (.Y(N448),.A(N401));
BUFX1 uut149 (.Y(N449),.A(N402));
BUFX1 uut150 (.Y(N450),.A(N403));
INVX1 uut151 (.Y(N451),.A(N424));
NOR2X1 uut152 (.Y(N460),.A(N406),.B(N425));
NOR2X1 uut153 (.Y(N463),.A(N409),.B(N426));
NAND2X1 uut154 (.Y(N466),.A(N442),.B(N410));
AND2X1 uut155 (.Y(N475),.A(N143fo0),.B(N427fo0));
AND2X1 uut156 (.Y(N476),.A(N310fo1),.B(N432fo0));
AND2X1 uut157 (.Y(N477),.A(N146fo0),.B(N427fo1));
AND2X1 uut158 (.Y(N478),.A(N310fo2),.B(N432fo1));
AND2X1 uut159 (.Y(N479),.A(N149fo0),.B(N427fo2));
AND2X1 uut160 (.Y(N480),.A(N310fo3),.B(N432fo2));
AND2X1 uut161 (.Y(N481),.A(N153fo0),.B(N427fo3));
AND2X1 uut162 (.Y(N482),.A(N310fo4),.B(N432fo3));
NAND2X1 uut163 (.Y(N483),.A(N443),.B(N1fo5));
OR2X1 uut164 (.Y(N488),.A(N369fo1),.B(N437fo0));
OR2X1 uut165 (.Y(N489),.A(N369fo2),.B(N437fo1));
OR2X1 uut166 (.Y(N490),.A(N369fo3),.B(N437fo2));
OR2X1 uut167 (.Y(N491),.A(N369fo4),.B(N437fo3));
NOR2X1 uut168 (.Y(N492),.A(N413),.B(N444));
NOR2X1 uut169 (.Y(N495),.A(N416),.B(N445));
NAND2X1 uut170 (.Y(N498),.A(N130fo0),.B(N460fo0));
OR2X1 uut171 (.Y(N499),.A(N130fo1),.B(N460fo1));
NAND2X1 uut172 (.Y(N500),.A(N463fo0),.B(N135fo0));
OR2X1 uut173 (.Y(N501),.A(N463fo1),.B(N135fo1));
AND2X1 uut174 (.Y(N502),.A(N91fo3),.B(N466fo0));
NOR2X1 uut175 (.Y(N503),.A(N475),.B(N476));
AND2X1 uut176 (.Y(N504),.A(N96fo3),.B(N466fo1));
NOR2X1 uut177 (.Y(N505),.A(N477),.B(N478));
AND2X1 uut178 (.Y(N506),.A(N101fo3),.B(N466fo2));
NOR2X1 uut179 (.Y(N507),.A(N479),.B(N480));
AND2X1 uut180 (.Y(N508),.A(N106fo3),.B(N466fo3));
NOR2X1 uut181 (.Y(N509),.A(N481),.B(N482));
AND2X1 uut182 (.Y(N510),.A(N143fo1),.B(N483fo0));
AND2X1 uut183 (.Y(N511),.A(N111fo3),.B(N466fo4));
AND2X1 uut184 (.Y(N512),.A(N146fo1),.B(N483fo1));
AND2X1 uut185 (.Y(N513),.A(N116fo3),.B(N466fo5));
AND2X1 uut186 (.Y(N514),.A(N149fo1),.B(N483fo2));
AND2X1 uut187 (.Y(N515),.A(N121fo3),.B(N466fo6));
AND2X1 uut188 (.Y(N516),.A(N153fo1),.B(N483fo3));
AND2X1 uut189 (.Y(N517),.A(N126fo2),.B(N466fo7));
NAND2X1 uut190 (.Y(N518),.A(N130fo2),.B(N492fo0));
OR2X1 uut191 (.Y(N519),.A(N130fo3),.B(N492fo1));
NAND2X1 uut192 (.Y(N520),.A(N495fo0),.B(N207fo0));
OR2X1 uut193 (.Y(N521),.A(N495fo1),.B(N207fo1));
AND2X1 uut194 (.Y(N522),.A(N451fo0),.B(N159fo2));
AND2X1 uut195 (.Y(N523),.A(N451fo1),.B(N165fo2));
AND2X1 uut196 (.Y(N524),.A(N451fo2),.B(N171fo2));
AND2X1 uut197 (.Y(N525),.A(N451fo3),.B(N177fo2));
AND2X1 uut198 (.Y(N526),.A(N451fo4),.B(N183fo2));
NAND2X1 uut199 (.Y(N527),.A(N451fo5),.B(N189fo2));
NAND2X1 uut200 (.Y(N528),.A(N451fo6),.B(N195fo2));
NAND2X1 uut201 (.Y(N529),.A(N451fo7),.B(N201fo2));
NAND2X1 uut202 (.Y(N530),.A(N498),.B(N499));
NAND2X1 uut203 (.Y(N533),.A(N500),.B(N501));
NOR2X1 uut204 (.Y(N536),.A(N309),.B(N502));
NOR2X1 uut205 (.Y(N537),.A(N316),.B(N504));
NOR2X1 uut206 (.Y(N538),.A(N317),.B(N506));
NOR2X1 uut207 (.Y(N539),.A(N318),.B(N508));
NOR2X1 uut208 (.Y(N540),.A(N510),.B(N511));
NOR2X1 uut209 (.Y(N541),.A(N512),.B(N513));
NOR2X1 uut210 (.Y(N542),.A(N514),.B(N515));
NOR2X1 uut211 (.Y(N543),.A(N516),.B(N517));
NAND2X1 uut212 (.Y(N544),.A(N518),.B(N519));
NAND2X1 uut213 (.Y(N547),.A(N520),.B(N521));
INVX1 uut214 (.Y(N550),.A(N530fo0));
INVX1 uut215 (.Y(N551),.A(N533fo0));
AND2X1 uut216 (.Y(N552),.A(N530fo1),.B(N533fo1));
NAND2X1 uut217 (.Y(N553),.A(N536),.B(N503));
NAND2X1 uut218 (.Y(N557),.A(N537),.B(N505));
NAND2X1 uut219 (.Y(N561),.A(N538),.B(N507));
NAND2X1 uut220 (.Y(N565),.A(N539),.B(N509));
NAND2X1 uut221 (.Y(N569),.A(N488),.B(N540));
NAND2X1 uut222 (.Y(N573),.A(N489),.B(N541));
NAND2X1 uut223 (.Y(N577),.A(N490),.B(N542));
NAND2X1 uut224 (.Y(N581),.A(N491),.B(N543));
INVX1 uut225 (.Y(N585),.A(N544fo0));
INVX1 uut226 (.Y(N586),.A(N547fo0));
AND2X1 uut227 (.Y(N587),.A(N544fo1),.B(N547fo1));
AND2X1 uut228 (.Y(N588),.A(N550),.B(N551));
AND2X1 uut229 (.Y(N589),.A(N585),.B(N586));
NAND2X1 uut230 (.Y(N590),.A(N553fo0),.B(N159fo3));
OR2X1 uut231 (.Y(N593),.A(N553fo1),.B(N159fo4));
AND2X1 uut232 (.Y(N596),.A(N246fo0),.B(N553fo2));
NAND2X1 uut233 (.Y(N597),.A(N557fo0),.B(N165fo3));
OR2X1 uut234 (.Y(N600),.A(N557fo1),.B(N165fo4));
AND2X1 uut235 (.Y(N605),.A(N246fo1),.B(N557fo2));
NAND2X1 uut236 (.Y(N606),.A(N561fo0),.B(N171fo3));
OR2X1 uut237 (.Y(N609),.A(N561fo1),.B(N171fo4));
AND2X1 uut238 (.Y(N615),.A(N246fo2),.B(N561fo2));
NAND2X1 uut239 (.Y(N616),.A(N565fo0),.B(N177fo3));
OR2X1 uut240 (.Y(N619),.A(N565fo1),.B(N177fo4));
AND2X1 uut241 (.Y(N624),.A(N246fo3),.B(N565fo2));
NAND2X1 uut242 (.Y(N625),.A(N569fo0),.B(N183fo3));
OR2X1 uut243 (.Y(N628),.A(N569fo1),.B(N183fo4));
AND2X1 uut244 (.Y(N631),.A(N246fo4),.B(N569fo2));
NAND2X1 uut245 (.Y(N632),.A(N573fo0),.B(N189fo3));
OR2X1 uut246 (.Y(N635),.A(N573fo1),.B(N189fo4));
AND2X1 uut247 (.Y(N640),.A(N246fo5),.B(N573fo2));
NAND2X1 uut248 (.Y(N641),.A(N577fo0),.B(N195fo3));
OR2X1 uut249 (.Y(N644),.A(N577fo1),.B(N195fo4));
AND2X1 uut250 (.Y(N650),.A(N246fo6),.B(N577fo2));
NAND2X1 uut251 (.Y(N651),.A(N581fo0),.B(N201fo3));
OR2X1 uut252 (.Y(N654),.A(N581fo1),.B(N201fo4));
AND2X1 uut253 (.Y(N659),.A(N246fo7),.B(N581fo2));
NOR2X1 uut254 (.Y(N660),.A(N552),.B(N588));
NOR2X1 uut255 (.Y(N661),.A(N587),.B(N589));
INVX1 uut256 (.Y(N662),.A(N590fo0));
AND2X1 uut257 (.Y(N665),.A(N593fo0),.B(N590fo1));
NOR2X1 uut258 (.Y(N669),.A(N596),.B(N522));
INVX1 uut259 (.Y(N670),.A(N597fo0));
AND2X1 uut260 (.Y(N673),.A(N600fo0),.B(N597fo1));
NOR2X1 uut261 (.Y(N677),.A(N605),.B(N523));
INVX1 uut262 (.Y(N678),.A(N606fo0));
AND2X1 uut263 (.Y(N682),.A(N609fo0),.B(N606fo1));
NOR2X1 uut264 (.Y(N686),.A(N615),.B(N524));
INVX1 uut265 (.Y(N687),.A(N616fo0));
AND2X1 uut266 (.Y(N692),.A(N619fo0),.B(N616fo1));
NOR2X1 uut267 (.Y(N696),.A(N624),.B(N525));
INVX1 uut268 (.Y(N697),.A(N625fo0));
AND2X1 uut269 (.Y(N700),.A(N628fo0),.B(N625fo1));
NOR2X1 uut270 (.Y(N704),.A(N631),.B(N526));
INVX1 uut271 (.Y(N705),.A(N632fo0));
AND2X1 uut272 (.Y(N708),.A(N635fo0),.B(N632fo1));
NOR2X1 uut273 (.Y(N712),.A(N337),.B(N640));
INVX1 uut274 (.Y(N713),.A(N641fo0));
AND2X1 uut275 (.Y(N717),.A(N644fo0),.B(N641fo1));
NOR2X1 uut276 (.Y(N721),.A(N339),.B(N650));
INVX1 uut277 (.Y(N722),.A(N651fo0));
AND2X1 uut278 (.Y(N727),.A(N654fo0),.B(N651fo1));
NOR2X1 uut279 (.Y(N731),.A(N341),.B(N659));
NAND2X1 uut280 (.Y(N732),.A(N654fo1),.B(N261fo0));
AND2X1 uut281 (.Y(ttmp49),.A(N654fo2),.B(N261fo1));
NAND2X1 uut282 (.Y(N733),.A(N644fo1),.B(ttmp49));
AND2X1 uut283 (.Y(ttmp51),.A(N654fo3),.B(N261fo2));
AND2X1 uut284 (.Y(ttmp52),.A(N635fo1),.B(ttmp51));
NAND2X1 uut285 (.Y(N734),.A(N644fo2),.B(ttmp52));
INVX1 uut286 (.Y(N735),.A(N662fo0));
AND2X1 uut287 (.Y(N736),.A(N228fo0),.B(N665fo0));
AND2X1 uut288 (.Y(N737),.A(N237fo0),.B(N662fo1));
INVX1 uut289 (.Y(N738),.A(N670fo0));
AND2X1 uut290 (.Y(N739),.A(N228fo1),.B(N673fo0));
AND2X1 uut291 (.Y(N740),.A(N237fo1),.B(N670fo1));
INVX1 uut292 (.Y(N741),.A(N678fo0));
AND2X1 uut293 (.Y(N742),.A(N228fo2),.B(N682fo0));
AND2X1 uut294 (.Y(N743),.A(N237fo2),.B(N678fo1));
INVX1 uut295 (.Y(N744),.A(N687fo0));
AND2X1 uut296 (.Y(N745),.A(N228fo3),.B(N692fo0));
AND2X1 uut297 (.Y(N746),.A(N237fo3),.B(N687fo1));
INVX1 uut298 (.Y(N747),.A(N697fo0));
AND2X1 uut299 (.Y(N748),.A(N228fo4),.B(N700fo0));
AND2X1 uut300 (.Y(N749),.A(N237fo4),.B(N697fo1));
INVX1 uut301 (.Y(N750),.A(N705fo0));
AND2X1 uut302 (.Y(N751),.A(N228fo5),.B(N708fo0));
AND2X1 uut303 (.Y(N752),.A(N237fo5),.B(N705fo1));
INVX1 uut304 (.Y(N753),.A(N713fo0));
AND2X1 uut305 (.Y(N754),.A(N228fo6),.B(N717fo0));
AND2X1 uut306 (.Y(N755),.A(N237fo6),.B(N713fo1));
INVX1 uut307 (.Y(N756),.A(N722fo0));
NOR2X1 uut308 (.Y(N757),.A(N727fo0),.B(N261fo3));
AND2X1 uut309 (.Y(N758),.A(N727fo1),.B(N261fo4));
AND2X1 uut310 (.Y(N759),.A(N228fo7),.B(N727fo2));
AND2X1 uut311 (.Y(N760),.A(N237fo7),.B(N722fo1));
NAND2X1 uut312 (.Y(N761),.A(N644fo3),.B(N722fo2));
NAND2X1 uut313 (.Y(N762),.A(N635fo2),.B(N713fo2));
AND2X1 uut314 (.Y(ttmp54),.A(N644fo4),.B(N722fo3));
NAND2X1 uut315 (.Y(N763),.A(N635fo3),.B(ttmp54));
NAND2X1 uut316 (.Y(N764),.A(N609fo1),.B(N687fo2));
NAND2X1 uut317 (.Y(N765),.A(N600fo1),.B(N678fo2));
AND2X1 uut318 (.Y(ttmp56),.A(N609fo2),.B(N687fo3));
NAND2X1 uut319 (.Y(N766),.A(N600fo2),.B(ttmp56));
BUFX1 uut320 (.Y(N767),.A(N660));
BUFX1 uut321 (.Y(N768),.A(N661));
NOR2X1 uut322 (.Y(N769),.A(N736),.B(N737));
NOR2X1 uut323 (.Y(N770),.A(N739),.B(N740));
NOR2X1 uut324 (.Y(N771),.A(N742),.B(N743));
NOR2X1 uut325 (.Y(N772),.A(N745),.B(N746));
AND2X1 uut326 (.Y(ttmp58),.A(N763),.B(N734));
AND2X1 uut327 (.Y(ttmp59),.A(N750),.B(ttmp58));
NAND2X1 uut328 (.Y(N773),.A(N762),.B(ttmp59));
NOR2X1 uut329 (.Y(N777),.A(N748),.B(N749));
AND2X1 uut330 (.Y(ttmp61),.A(N761),.B(N733));
NAND2X1 uut331 (.Y(N778),.A(N753),.B(ttmp61));
NOR2X1 uut332 (.Y(N781),.A(N751),.B(N752));
NAND2X1 uut333 (.Y(N782),.A(N756),.B(N732));
NOR2X1 uut334 (.Y(N785),.A(N754),.B(N755));
NOR2X1 uut335 (.Y(N786),.A(N757),.B(N758));
NOR2X1 uut336 (.Y(N787),.A(N759),.B(N760));
NOR2X1 uut337 (.Y(N788),.A(N700fo1),.B(N773fo0));
AND2X1 uut338 (.Y(N789),.A(N700fo2),.B(N773fo1));
NOR2X1 uut339 (.Y(N790),.A(N708fo1),.B(N778fo0));
AND2X1 uut340 (.Y(N791),.A(N708fo2),.B(N778fo1));
NOR2X1 uut341 (.Y(N792),.A(N717fo1),.B(N782fo0));
AND2X1 uut342 (.Y(N793),.A(N717fo2),.B(N782fo1));
AND2X1 uut343 (.Y(N794),.A(N219fo0),.B(N786));
NAND2X1 uut344 (.Y(N795),.A(N628fo1),.B(N773fo2));
NAND2X1 uut345 (.Y(N796),.A(N795),.B(N747));
NOR2X1 uut346 (.Y(N802),.A(N788),.B(N789));
NOR2X1 uut347 (.Y(N803),.A(N790),.B(N791));
NOR2X1 uut348 (.Y(N804),.A(N792),.B(N793));
NOR2X1 uut349 (.Y(N805),.A(N340),.B(N794));
NOR2X1 uut350 (.Y(N806),.A(N692fo1),.B(N796fo0));
AND2X1 uut351 (.Y(N807),.A(N692fo2),.B(N796fo1));
AND2X1 uut352 (.Y(N808),.A(N219fo1),.B(N802));
AND2X1 uut353 (.Y(N809),.A(N219fo2),.B(N803));
AND2X1 uut354 (.Y(N810),.A(N219fo3),.B(N804));
AND2X1 uut355 (.Y(ttmp63),.A(N731),.B(N529));
AND2X1 uut356 (.Y(ttmp64),.A(N805),.B(ttmp63));
NAND2X1 uut357 (.Y(N811),.A(N787),.B(ttmp64));
NAND2X1 uut358 (.Y(N812),.A(N619fo1),.B(N796fo2));
AND2X1 uut359 (.Y(ttmp66),.A(N619fo2),.B(N796fo3));
NAND2X1 uut360 (.Y(N813),.A(N609fo3),.B(ttmp66));
AND2X1 uut361 (.Y(ttmp68),.A(N619fo3),.B(N796fo4));
AND2X1 uut362 (.Y(ttmp69),.A(N600fo3),.B(ttmp68));
NAND2X1 uut363 (.Y(N814),.A(N609fo4),.B(ttmp69));
AND2X1 uut364 (.Y(ttmp71),.A(N766),.B(N814));
AND2X1 uut365 (.Y(ttmp72),.A(N738),.B(ttmp71));
NAND2X1 uut366 (.Y(N815),.A(N765),.B(ttmp72));
AND2X1 uut367 (.Y(ttmp74),.A(N764),.B(N813));
NAND2X1 uut368 (.Y(N819),.A(N741),.B(ttmp74));
NAND2X1 uut369 (.Y(N822),.A(N744),.B(N812));
NOR2X1 uut370 (.Y(N825),.A(N806),.B(N807));
NOR2X1 uut371 (.Y(N826),.A(N335),.B(N808));
NOR2X1 uut372 (.Y(N827),.A(N336),.B(N809));
NOR2X1 uut373 (.Y(N828),.A(N338),.B(N810));
INVX1 uut374 (.Y(N829),.A(N811));
NOR2X1 uut375 (.Y(N830),.A(N665fo1),.B(N815fo0));
AND2X1 uut376 (.Y(N831),.A(N665fo2),.B(N815fo1));
NOR2X1 uut377 (.Y(N832),.A(N673fo1),.B(N819fo0));
AND2X1 uut378 (.Y(N833),.A(N673fo2),.B(N819fo1));
NOR2X1 uut379 (.Y(N834),.A(N682fo1),.B(N822fo0));
AND2X1 uut380 (.Y(N835),.A(N682fo2),.B(N822fo1));
AND2X1 uut381 (.Y(N836),.A(N219fo4),.B(N825));
AND2X1 uut382 (.Y(ttmp76),.A(N777),.B(N704));
NAND2X1 uut383 (.Y(N837),.A(N826),.B(ttmp76));
AND2X1 uut384 (.Y(ttmp78),.A(N712),.B(N527));
AND2X1 uut385 (.Y(ttmp79),.A(N827),.B(ttmp78));
NAND2X1 uut386 (.Y(N838),.A(N781),.B(ttmp79));
AND2X1 uut387 (.Y(ttmp81),.A(N721),.B(N528));
AND2X1 uut388 (.Y(ttmp82),.A(N828),.B(ttmp81));
NAND2X1 uut389 (.Y(N839),.A(N785),.B(ttmp82));
INVX1 uut390 (.Y(N840),.A(N829));
NAND2X1 uut391 (.Y(N841),.A(N815fo2),.B(N593fo1));
NOR2X1 uut392 (.Y(N842),.A(N830),.B(N831));
NOR2X1 uut393 (.Y(N843),.A(N832),.B(N833));
NOR2X1 uut394 (.Y(N844),.A(N834),.B(N835));
NOR2X1 uut395 (.Y(N845),.A(N334),.B(N836));
INVX1 uut396 (.Y(N846),.A(N837));
INVX1 uut397 (.Y(N847),.A(N838));
INVX1 uut398 (.Y(N848),.A(N839));
AND2X1 uut399 (.Y(N849),.A(N735),.B(N841));
BUFX1 uut400 (.Y(N850),.A(N840));
AND2X1 uut401 (.Y(N851),.A(N219fo5),.B(N842));
AND2X1 uut402 (.Y(N852),.A(N219fo6),.B(N843));
AND2X1 uut403 (.Y(N853),.A(N219fo7),.B(N844));
AND2X1 uut404 (.Y(ttmp84),.A(N772),.B(N696));
NAND2X1 uut405 (.Y(N854),.A(N845),.B(ttmp84));
INVX1 uut406 (.Y(N855),.A(N846));
INVX1 uut407 (.Y(N856),.A(N847));
INVX1 uut408 (.Y(N857),.A(N848));
INVX1 uut409 (.Y(N858),.A(N849));
NOR2X1 uut410 (.Y(N859),.A(N417),.B(N851));
NOR2X1 uut411 (.Y(N860),.A(N332),.B(N852));
NOR2X1 uut412 (.Y(N861),.A(N333),.B(N853));
INVX1 uut413 (.Y(N862),.A(N854));
BUFX1 uut414 (.Y(N863),.A(N855));
BUFX1 uut415 (.Y(N864),.A(N856));
BUFX1 uut416 (.Y(N865),.A(N857));
BUFX1 uut417 (.Y(N866),.A(N858));
AND2X1 uut418 (.Y(ttmp86),.A(N769),.B(N669));
NAND2X1 uut419 (.Y(N867),.A(N859),.B(ttmp86));
AND2X1 uut420 (.Y(ttmp88),.A(N770),.B(N677));
NAND2X1 uut421 (.Y(N868),.A(N860),.B(ttmp88));
AND2X1 uut422 (.Y(ttmp90),.A(N771),.B(N686));
NAND2X1 uut423 (.Y(N869),.A(N861),.B(ttmp90));
INVX1 uut424 (.Y(N870),.A(N862));
INVX1 uut425 (.Y(N871),.A(N867));
INVX1 uut426 (.Y(N872),.A(N868));
INVX1 uut427 (.Y(N873),.A(N869));
BUFX1 uut428 (.Y(N874),.A(N870));
INVX1 uut429 (.Y(N875),.A(N871));
INVX1 uut430 (.Y(N876),.A(N872));
INVX1 uut431 (.Y(N877),.A(N873));
BUFX1 uut432 (.Y(N878),.A(N875));
BUFX1 uut433 (.Y(N879),.A(N876));
BUFX1 uut434 (.Y(N880),.A(N877));
fanout6 uut_fo0 (.A(N1),.Y1(N1fo0),.Y2(N1fo1),.Y3(N1fo2),.Y4(N1fo3),.Y5(N1fo4),.Y6(N1fo5));
fanout4 uut_fo1 (.A(N8),.Y1(N8fo0),.Y2(N8fo1),.Y3(N8fo2),.Y4(N8fo3));
fanout3 uut_fo2 (.A(N13),.Y1(N13fo0),.Y2(N13fo1),.Y3(N13fo2));
fanout8 uut_fo3 (.A(N17),.Y1(N17fo0),.Y2(N17fo1),.Y3(N17fo2),.Y4(N17fo3),.Y5(N17fo4),.Y6(N17fo5),.Y7(N17fo6),.Y8(N17fo7));
fanout2 uut_fo4 (.A(N26),.Y1(N26fo0),.Y2(N26fo1));
fanout6 uut_fo5 (.A(N29),.Y1(N29fo0),.Y2(N29fo1),.Y3(N29fo2),.Y4(N29fo3),.Y5(N29fo4),.Y6(N29fo5));
fanout5 uut_fo6 (.A(N36),.Y1(N36fo0),.Y2(N36fo1),.Y3(N36fo2),.Y4(N36fo3),.Y5(N36fo4));
fanout8 uut_fo7 (.A(N42),.Y1(N42fo0),.Y2(N42fo1),.Y3(N42fo2),.Y4(N42fo3),.Y5(N42fo4),.Y6(N42fo5),.Y7(N42fo6),.Y8(N42fo7));
fanout3 uut_fo8 (.A(N51),.Y1(N51fo0),.Y2(N51fo1),.Y3(N51fo2));
fanout3 uut_fo9 (.A(N55),.Y1(N55fo0),.Y2(N55fo1),.Y3(N55fo2));
fanout8 uut_fo10 (.A(N59),.Y1(N59fo0),.Y2(N59fo1),.Y3(N59fo2),.Y4(N59fo3),.Y5(N59fo4),.Y6(N59fo5),.Y7(N59fo6),.Y8(N59fo7));
fanout3 uut_fo11 (.A(N68),.Y1(N68fo0),.Y2(N68fo1),.Y3(N68fo2));
fanout4 uut_fo15 (.A(N75),.Y1(N75fo0),.Y2(N75fo1),.Y3(N75fo2),.Y4(N75fo3));
fanout4 uut_fo16 (.A(N80),.Y1(N80fo0),.Y2(N80fo1),.Y3(N80fo2),.Y4(N80fo3));
fanout4 uut_fo23 (.A(N91),.Y1(N91fo0),.Y2(N91fo1),.Y3(N91fo2),.Y4(N91fo3));
fanout4 uut_fo24 (.A(N96),.Y1(N96fo0),.Y2(N96fo1),.Y3(N96fo2),.Y4(N96fo3));
fanout4 uut_fo25 (.A(N101),.Y1(N101fo0),.Y2(N101fo1),.Y3(N101fo2),.Y4(N101fo3));
fanout4 uut_fo26 (.A(N106),.Y1(N106fo0),.Y2(N106fo1),.Y3(N106fo2),.Y4(N106fo3));
fanout4 uut_fo27 (.A(N111),.Y1(N111fo0),.Y2(N111fo1),.Y3(N111fo2),.Y4(N111fo3));
fanout4 uut_fo28 (.A(N116),.Y1(N116fo0),.Y2(N116fo1),.Y3(N116fo2),.Y4(N116fo3));
fanout4 uut_fo29 (.A(N121),.Y1(N121fo0),.Y2(N121fo1),.Y3(N121fo2),.Y4(N121fo3));
fanout3 uut_fo30 (.A(N126),.Y1(N126fo0),.Y2(N126fo1),.Y3(N126fo2));
fanout4 uut_fo31 (.A(N130),.Y1(N130fo0),.Y2(N130fo1),.Y3(N130fo2),.Y4(N130fo3));
fanout2 uut_fo32 (.A(N135),.Y1(N135fo0),.Y2(N135fo1));
fanout4 uut_fo33 (.A(N138),.Y1(N138fo0),.Y2(N138fo1),.Y3(N138fo2),.Y4(N138fo3));
fanout2 uut_fo34 (.A(N143),.Y1(N143fo0),.Y2(N143fo1));
fanout2 uut_fo35 (.A(N146),.Y1(N146fo0),.Y2(N146fo1));
fanout2 uut_fo36 (.A(N149),.Y1(N149fo0),.Y2(N149fo1));
fanout2 uut_fo38 (.A(N153),.Y1(N153fo0),.Y2(N153fo1));
fanout2 uut_fo39 (.A(N156),.Y1(N156fo0),.Y2(N156fo1));
fanout5 uut_fo40 (.A(N159),.Y1(N159fo0),.Y2(N159fo1),.Y3(N159fo2),.Y4(N159fo3),.Y5(N159fo4));
fanout5 uut_fo41 (.A(N165),.Y1(N165fo0),.Y2(N165fo1),.Y3(N165fo2),.Y4(N165fo3),.Y5(N165fo4));
fanout5 uut_fo42 (.A(N171),.Y1(N171fo0),.Y2(N171fo1),.Y3(N171fo2),.Y4(N171fo3),.Y5(N171fo4));
fanout5 uut_fo43 (.A(N177),.Y1(N177fo0),.Y2(N177fo1),.Y3(N177fo2),.Y4(N177fo3),.Y5(N177fo4));
fanout5 uut_fo44 (.A(N183),.Y1(N183fo0),.Y2(N183fo1),.Y3(N183fo2),.Y4(N183fo3),.Y5(N183fo4));
fanout5 uut_fo45 (.A(N189),.Y1(N189fo0),.Y2(N189fo1),.Y3(N189fo2),.Y4(N189fo3),.Y5(N189fo4));
fanout5 uut_fo46 (.A(N195),.Y1(N195fo0),.Y2(N195fo1),.Y3(N195fo2),.Y4(N195fo3),.Y5(N195fo4));
fanout5 uut_fo47 (.A(N201),.Y1(N201fo0),.Y2(N201fo1),.Y3(N201fo2),.Y4(N201fo3),.Y5(N201fo4));
fanout2 uut_fo48 (.A(N207),.Y1(N207fo0),.Y2(N207fo1));
fanout8 uut_fo49 (.A(N210),.Y1(N210fo0),.Y2(N210fo1),.Y3(N210fo2),.Y4(N210fo3),.Y5(N210fo4),.Y6(N210fo5),.Y7(N210fo6),.Y8(N210fo7));
fanout8 uut_fo50 (.A(N219),.Y1(N219fo0),.Y2(N219fo1),.Y3(N219fo2),.Y4(N219fo3),.Y5(N219fo4),.Y6(N219fo5),.Y7(N219fo6),.Y8(N219fo7));
fanout8 uut_fo51 (.A(N228),.Y1(N228fo0),.Y2(N228fo1),.Y3(N228fo2),.Y4(N228fo3),.Y5(N228fo4),.Y6(N228fo5),.Y7(N228fo6),.Y8(N228fo7));
fanout8 uut_fo52 (.A(N237),.Y1(N237fo0),.Y2(N237fo1),.Y3(N237fo2),.Y4(N237fo3),.Y5(N237fo4),.Y6(N237fo5),.Y7(N237fo6),.Y8(N237fo7));
fanout8 uut_fo53 (.A(N246),.Y1(N246fo0),.Y2(N246fo1),.Y3(N246fo2),.Y4(N246fo3),.Y5(N246fo4),.Y6(N246fo5),.Y7(N246fo6),.Y8(N246fo7));
fanout3 uut_fo54 (.A(N255),.Y1(N255fo0),.Y2(N255fo1),.Y3(N255fo2));
fanout5 uut_fo57 (.A(N261),.Y1(N261fo0),.Y2(N261fo1),.Y3(N261fo2),.Y4(N261fo3),.Y5(N261fo4));
fanout2 uut_fo_w1 (.A(N606),.Y1(N606fo0),.Y2(N606fo1));
fanout2 uut_fo_w2 (.A(N544),.Y1(N544fo0),.Y2(N544fo1));
fanout2 uut_fo_w3 (.A(N593),.Y1(N593fo0),.Y2(N593fo1));
fanout3 uut_fo_w13 (.A(N553),.Y1(N553fo0),.Y2(N553fo1),.Y3(N553fo2));
fanout2 uut_fo_w14 (.A(N460),.Y1(N460fo0),.Y2(N460fo1));
fanout3 uut_fo_w48 (.A(N665),.Y1(N665fo0),.Y2(N665fo1),.Y3(N665fo2));
fanout2 uut_fo_w58 (.A(N287),.Y1(N287fo0),.Y2(N287fo1));
fanout5 uut_fo_w68 (.A(N369),.Y1(N369fo0),.Y2(N369fo1),.Y3(N369fo2),.Y4(N369fo3),.Y5(N369fo4));
fanout2 uut_fo_w74 (.A(N782),.Y1(N782fo0),.Y2(N782fo1));
fanout2 uut_fo_w82 (.A(N463),.Y1(N463fo0),.Y2(N463fo1));
fanout2 uut_fo_w87 (.A(N382),.Y1(N382fo0),.Y2(N382fo1));
fanout3 uut_fo_w88 (.A(N565),.Y1(N565fo0),.Y2(N565fo1),.Y3(N565fo2));
fanout3 uut_fo_w91 (.A(N682),.Y1(N682fo0),.Y2(N682fo1),.Y3(N682fo2));
fanout5 uut_fo_w92 (.A(N796),.Y1(N796fo0),.Y2(N796fo1),.Y3(N796fo2),.Y4(N796fo3),.Y5(N796fo4));
fanout2 uut_fo_w94 (.A(N819),.Y1(N819fo0),.Y2(N819fo1));
fanout5 uut_fo_w99 (.A(N310),.Y1(N310fo0),.Y2(N310fo1),.Y3(N310fo2),.Y4(N310fo3),.Y5(N310fo4));
fanout2 uut_fo_w100 (.A(N597),.Y1(N597fo0),.Y2(N597fo1));
fanout2 uut_fo_w101 (.A(N385),.Y1(N385fo0),.Y2(N385fo1));
fanout3 uut_fo_w110 (.A(N581),.Y1(N581fo0),.Y2(N581fo1),.Y3(N581fo2));
fanout2 uut_fo_w111 (.A(N625),.Y1(N625fo0),.Y2(N625fo1));
fanout3 uut_fo_w124 (.A(N815),.Y1(N815fo0),.Y2(N815fo1),.Y3(N815fo2));
fanout2 uut_fo_w132 (.A(N590),.Y1(N590fo0),.Y2(N590fo1));
fanout3 uut_fo_w135 (.A(N700),.Y1(N700fo0),.Y2(N700fo1),.Y3(N700fo2));
fanout3 uut_fo_w139 (.A(N692),.Y1(N692fo0),.Y2(N692fo1),.Y3(N692fo2));
fanout5 uut_fo_w145 (.A(N609),.Y1(N609fo0),.Y2(N609fo1),.Y3(N609fo2),.Y4(N609fo3),.Y5(N609fo4));
fanout3 uut_fo_w146 (.A(N773),.Y1(N773fo0),.Y2(N773fo1),.Y3(N773fo2));
fanout2 uut_fo_w150 (.A(N270),.Y1(N270fo0),.Y2(N270fo1));
fanout2 uut_fo_w151 (.A(N366),.Y1(N366fo0),.Y2(N366fo1));
fanout3 uut_fo_w157 (.A(N713),.Y1(N713fo0),.Y2(N713fo1),.Y3(N713fo2));
fanout2 uut_fo_w165 (.A(N778),.Y1(N778fo0),.Y2(N778fo1));
fanout3 uut_fo_w175 (.A(N280),.Y1(N280fo0),.Y2(N280fo1),.Y3(N280fo2));
fanout3 uut_fo_w177 (.A(N573),.Y1(N573fo0),.Y2(N573fo1),.Y3(N573fo2));
fanout2 uut_fo_w179 (.A(N628),.Y1(N628fo0),.Y2(N628fo1));
fanout3 uut_fo_w186 (.A(N708),.Y1(N708fo0),.Y2(N708fo1),.Y3(N708fo2));
fanout4 uut_fo_w190 (.A(N437),.Y1(N437fo0),.Y2(N437fo1),.Y3(N437fo2),.Y4(N437fo3));
fanout2 uut_fo_w203 (.A(N547),.Y1(N547fo0),.Y2(N547fo1));
fanout2 uut_fo_w208 (.A(N276),.Y1(N276fo0),.Y2(N276fo1));
fanout2 uut_fo_w217 (.A(N492),.Y1(N492fo0),.Y2(N492fo1));
fanout2 uut_fo_w222 (.A(N376),.Y1(N376fo0),.Y2(N376fo1));
fanout3 uut_fo_w235 (.A(N577),.Y1(N577fo0),.Y2(N577fo1),.Y3(N577fo2));
fanout2 uut_fo_w236 (.A(N357),.Y1(N357fo0),.Y2(N357fo1));
fanout4 uut_fo_w239 (.A(N654),.Y1(N654fo0),.Y2(N654fo1),.Y3(N654fo2),.Y4(N654fo3));
fanout4 uut_fo_w243 (.A(N687),.Y1(N687fo0),.Y2(N687fo1),.Y3(N687fo2),.Y4(N687fo3));
fanout3 uut_fo_w256 (.A(N717),.Y1(N717fo0),.Y2(N717fo1),.Y3(N717fo2));
fanout2 uut_fo_w258 (.A(N641),.Y1(N641fo0),.Y2(N641fo1));
fanout4 uut_fo_w259 (.A(N722),.Y1(N722fo0),.Y2(N722fo1),.Y3(N722fo2),.Y4(N722fo3));
fanout2 uut_fo_w260 (.A(N363),.Y1(N363fo0),.Y2(N363fo1));
fanout4 uut_fo_w261 (.A(N483),.Y1(N483fo0),.Y2(N483fo1),.Y3(N483fo2),.Y4(N483fo3));
fanout3 uut_fo_w264 (.A(N727),.Y1(N727fo0),.Y2(N727fo1),.Y3(N727fo2));
fanout3 uut_fo_w271 (.A(N678),.Y1(N678fo0),.Y2(N678fo1),.Y3(N678fo2));
fanout3 uut_fo_w273 (.A(N673),.Y1(N673fo0),.Y2(N673fo1),.Y3(N673fo2));
fanout4 uut_fo_w275 (.A(N432),.Y1(N432fo0),.Y2(N432fo1),.Y3(N432fo2),.Y4(N432fo3));
fanout2 uut_fo_w281 (.A(N273),.Y1(N273fo0),.Y2(N273fo1));
fanout2 uut_fo_w283 (.A(N697),.Y1(N697fo0),.Y2(N697fo1));
fanout5 uut_fo_w284 (.A(N393),.Y1(N393fo0),.Y2(N393fo1),.Y3(N393fo2),.Y4(N393fo3),.Y5(N393fo4));
fanout2 uut_fo_w290 (.A(N379),.Y1(N379fo0),.Y2(N379fo1));
fanout5 uut_fo_w292 (.A(N644),.Y1(N644fo0),.Y2(N644fo1),.Y3(N644fo2),.Y4(N644fo3),.Y5(N644fo4));
fanout4 uut_fo_w301 (.A(N427),.Y1(N427fo0),.Y2(N427fo1),.Y3(N427fo2),.Y4(N427fo3));
fanout2 uut_fo_w303 (.A(N298),.Y1(N298fo0),.Y2(N298fo1));
fanout2 uut_fo_w310 (.A(N670),.Y1(N670fo0),.Y2(N670fo1));
fanout2 uut_fo_w311 (.A(N495),.Y1(N495fo0),.Y2(N495fo1));
fanout2 uut_fo_w313 (.A(N360),.Y1(N360fo0),.Y2(N360fo1));
fanout2 uut_fo_w314 (.A(N822),.Y1(N822fo0),.Y2(N822fo1));
fanout2 uut_fo_w324 (.A(N651),.Y1(N651fo0),.Y2(N651fo1));
fanout8 uut_fo_w338 (.A(N466),.Y1(N466fo0),.Y2(N466fo1),.Y3(N466fo2),.Y4(N466fo3),.Y5(N466fo4),.Y6(N466fo5),.Y7(N466fo6),.Y8(N466fo7));
fanout3 uut_fo_w345 (.A(N561),.Y1(N561fo0),.Y2(N561fo1),.Y3(N561fo2));
fanout8 uut_fo_w353 (.A(N451),.Y1(N451fo0),.Y2(N451fo1),.Y3(N451fo2),.Y4(N451fo3),.Y5(N451fo4),.Y6(N451fo5),.Y7(N451fo6),.Y8(N451fo7));
fanout2 uut_fo_w363 (.A(N530),.Y1(N530fo0),.Y2(N530fo1));
fanout4 uut_fo_w365 (.A(N635),.Y1(N635fo0),.Y2(N635fo1),.Y3(N635fo2),.Y4(N635fo3));
fanout2 uut_fo_w366 (.A(N632),.Y1(N632fo0),.Y2(N632fo1));
fanout4 uut_fo_w370 (.A(N619),.Y1(N619fo0),.Y2(N619fo1),.Y3(N619fo2),.Y4(N619fo3));
fanout2 uut_fo_w373 (.A(N705),.Y1(N705fo0),.Y2(N705fo1));
fanout4 uut_fo_w375 (.A(N600),.Y1(N600fo0),.Y2(N600fo1),.Y3(N600fo2),.Y4(N600fo3));
fanout3 uut_fo_w376 (.A(N557),.Y1(N557fo0),.Y2(N557fo1),.Y3(N557fo2));
fanout3 uut_fo_w382 (.A(N569),.Y1(N569fo0),.Y2(N569fo1),.Y3(N569fo2));
fanout2 uut_fo_w385 (.A(N319),.Y1(N319fo0),.Y2(N319fo1));
fanout2 uut_fo_w386 (.A(N616),.Y1(N616fo0),.Y2(N616fo1));
fanout2 uut_fo_w405 (.A(N662),.Y1(N662fo0),.Y2(N662fo1));
fanout2 uut_fo_w407 (.A(N533),.Y1(N533fo0),.Y2(N533fo1));
endmodule
