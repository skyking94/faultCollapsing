module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,N137;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N1fo0,N5fo0,N9fo0,N13fo0,N17fo0,N21fo0,N25fo0,N29fo0,N33fo0,N37fo0,N41fo0,N45fo0,N49fo0,N53fo0,N57fo0,N61fo0,N65fo0,N69fo0,N73fo0,N77fo0,N81fo0,N85fo0,N89fo0,N93fo0,N97fo0,N101fo0,N105fo0,N109fo0,N113fo0,N117fo0,N121fo0,N125fo0,N137fo0,N137fo1,N137fo2,N137fo3,N137fo4,N137fo5,N137fo6,N137fo7,N1fo1,N17fo1,N33fo1,N49fo1,N5fo1,N21fo1,N37fo1,N53fo1,N9fo1,N25fo1,N41fo1,N57fo1,N13fo1,N29fo1,N45fo1,N61fo1,N65fo1,N81fo1,N97fo1,N113fo1,N69fo1,N85fo1,N101fo1,N117fo1,N73fo1,N89fo1,N105fo1,N121fo1,N77fo1,N93fo1,N109fo1,N125fo1,N290fo0,N293fo0,N296fo0,N299fo0,N290fo1,N296fo1,N293fo1,N299fo1,N302fo0,N305fo0,N308fo0,N311fo0,N302fo1,N308fo1,N305fo1,N311fo1,N354fo0,N367fo0,N380fo0,N354fo1,N367fo1,N393fo0,N354fo2,N380fo1,N393fo1,N367fo2,N380fo2,N393fo2,N419fo0,N445fo0,N419fo1,N432fo0,N406fo0,N445fo1,N406fo1,N432fo1,N406fo2,N419fo2,N432fo2,N406fo3,N419fo3,N445fo2,N406fo4,N432fo3,N445fo3,N419fo4,N432fo4,N445fo4,N367fo3,N393fo3,N367fo4,N380fo3,N354fo3,N393fo4,N354fo4,N380fo4,N393fo5,N380fo5,N367fo5,N354fo5,N445fo5,N432fo5,N419fo5,N406fo5,N602fo0,N406fo6,N432fo6,N445fo6,N602fo1,N406fo7,N602fo2,N419fo6,N432fo7,N445fo7,N602fo3,N419fo7,N607fo0,N354fo6,N380fo6,N393fo6,N607fo1,N354fo7,N607fo2,N367fo6,N380fo7,N393fo7,N607fo3,N367fo7,N354fo8,N620fo0,N367fo8,N620fo1,N380fo8,N620fo2,N393fo8,N620fo3,N354fo9,N625fo0,N367fo9,N625fo1,N380fo9,N625fo2,N393fo9,N625fo3,N354fo10,N630fo0,N367fo10,N630fo1,N380fo10,N630fo2,N393fo10,N630fo3,N354fo11,N635fo0,N367fo11,N635fo1,N380fo11,N635fo2,N393fo11,N635fo3,N406fo8,N640fo0,N419fo8,N640fo1,N432fo8,N640fo2,N445fo8,N640fo3,N406fo9,N645fo0,N419fo9,N645fo1,N432fo9,N645fo2,N445fo9,N645fo3,N406fo10,N650fo0,N419fo10,N650fo1,N432fo10,N650fo2,N445fo10,N650fo3,N406fo11,N655fo0,N419fo11,N655fo1,N432fo11,N655fo2,N445fo11,N655fo3,N1fo2,N5fo2,N9fo2,N13fo2,N17fo2,N21fo2,N25fo2,N29fo2,N33fo2,N37fo2,N41fo2,N45fo2,N49fo2,N53fo2,N57fo2,N61fo2,N65fo2,N69fo2,N73fo2,N77fo2,N81fo2,N85fo2,N89fo2,N93fo2,N97fo2,N101fo2,N105fo2,N109fo2,N113fo2,N117fo2,N121fo2,N125fo2;
XOR2X1 uut0 (.Y(N250),.A(N1fo0),.B(N5fo0));
XOR2X1 uut1 (.Y(N251),.A(N9fo0),.B(N13fo0));
XOR2X1 uut2 (.Y(N252),.A(N17fo0),.B(N21fo0));
XOR2X1 uut3 (.Y(N253),.A(N25fo0),.B(N29fo0));
XOR2X1 uut4 (.Y(N254),.A(N33fo0),.B(N37fo0));
XOR2X1 uut5 (.Y(N255),.A(N41fo0),.B(N45fo0));
XOR2X1 uut6 (.Y(N256),.A(N49fo0),.B(N53fo0));
XOR2X1 uut7 (.Y(N257),.A(N57fo0),.B(N61fo0));
XOR2X1 uut8 (.Y(N258),.A(N65fo0),.B(N69fo0));
XOR2X1 uut9 (.Y(N259),.A(N73fo0),.B(N77fo0));
XOR2X1 uut10 (.Y(N260),.A(N81fo0),.B(N85fo0));
XOR2X1 uut11 (.Y(N261),.A(N89fo0),.B(N93fo0));
XOR2X1 uut12 (.Y(N262),.A(N97fo0),.B(N101fo0));
XOR2X1 uut13 (.Y(N263),.A(N105fo0),.B(N109fo0));
XOR2X1 uut14 (.Y(N264),.A(N113fo0),.B(N117fo0));
XOR2X1 uut15 (.Y(N265),.A(N121fo0),.B(N125fo0));
AND2X1 uut16 (.Y(N266),.A(N129),.B(N137fo0));
AND2X1 uut17 (.Y(N267),.A(N130),.B(N137fo1));
AND2X1 uut18 (.Y(N268),.A(N131),.B(N137fo2));
AND2X1 uut19 (.Y(N269),.A(N132),.B(N137fo3));
AND2X1 uut20 (.Y(N270),.A(N133),.B(N137fo4));
AND2X1 uut21 (.Y(N271),.A(N134),.B(N137fo5));
AND2X1 uut22 (.Y(N272),.A(N135),.B(N137fo6));
AND2X1 uut23 (.Y(N273),.A(N136),.B(N137fo7));
XOR2X1 uut24 (.Y(N274),.A(N1fo1),.B(N17fo1));
XOR2X1 uut25 (.Y(N275),.A(N33fo1),.B(N49fo1));
XOR2X1 uut26 (.Y(N276),.A(N5fo1),.B(N21fo1));
XOR2X1 uut27 (.Y(N277),.A(N37fo1),.B(N53fo1));
XOR2X1 uut28 (.Y(N278),.A(N9fo1),.B(N25fo1));
XOR2X1 uut29 (.Y(N279),.A(N41fo1),.B(N57fo1));
XOR2X1 uut30 (.Y(N280),.A(N13fo1),.B(N29fo1));
XOR2X1 uut31 (.Y(N281),.A(N45fo1),.B(N61fo1));
XOR2X1 uut32 (.Y(N282),.A(N65fo1),.B(N81fo1));
XOR2X1 uut33 (.Y(N283),.A(N97fo1),.B(N113fo1));
XOR2X1 uut34 (.Y(N284),.A(N69fo1),.B(N85fo1));
XOR2X1 uut35 (.Y(N285),.A(N101fo1),.B(N117fo1));
XOR2X1 uut36 (.Y(N286),.A(N73fo1),.B(N89fo1));
XOR2X1 uut37 (.Y(N287),.A(N105fo1),.B(N121fo1));
XOR2X1 uut38 (.Y(N288),.A(N77fo1),.B(N93fo1));
XOR2X1 uut39 (.Y(N289),.A(N109fo1),.B(N125fo1));
XOR2X1 uut40 (.Y(N290),.A(N250),.B(N251));
XOR2X1 uut41 (.Y(N293),.A(N252),.B(N253));
XOR2X1 uut42 (.Y(N296),.A(N254),.B(N255));
XOR2X1 uut43 (.Y(N299),.A(N256),.B(N257));
XOR2X1 uut44 (.Y(N302),.A(N258),.B(N259));
XOR2X1 uut45 (.Y(N305),.A(N260),.B(N261));
XOR2X1 uut46 (.Y(N308),.A(N262),.B(N263));
XOR2X1 uut47 (.Y(N311),.A(N264),.B(N265));
XOR2X1 uut48 (.Y(N314),.A(N274),.B(N275));
XOR2X1 uut49 (.Y(N315),.A(N276),.B(N277));
XOR2X1 uut50 (.Y(N316),.A(N278),.B(N279));
XOR2X1 uut51 (.Y(N317),.A(N280),.B(N281));
XOR2X1 uut52 (.Y(N318),.A(N282),.B(N283));
XOR2X1 uut53 (.Y(N319),.A(N284),.B(N285));
XOR2X1 uut54 (.Y(N320),.A(N286),.B(N287));
XOR2X1 uut55 (.Y(N321),.A(N288),.B(N289));
XOR2X1 uut56 (.Y(N338),.A(N290fo0),.B(N293fo0));
XOR2X1 uut57 (.Y(N339),.A(N296fo0),.B(N299fo0));
XOR2X1 uut58 (.Y(N340),.A(N290fo1),.B(N296fo1));
XOR2X1 uut59 (.Y(N341),.A(N293fo1),.B(N299fo1));
XOR2X1 uut60 (.Y(N342),.A(N302fo0),.B(N305fo0));
XOR2X1 uut61 (.Y(N343),.A(N308fo0),.B(N311fo0));
XOR2X1 uut62 (.Y(N344),.A(N302fo1),.B(N308fo1));
XOR2X1 uut63 (.Y(N345),.A(N305fo1),.B(N311fo1));
XOR2X1 uut64 (.Y(N346),.A(N266),.B(N342));
XOR2X1 uut65 (.Y(N347),.A(N267),.B(N343));
XOR2X1 uut66 (.Y(N348),.A(N268),.B(N344));
XOR2X1 uut67 (.Y(N349),.A(N269),.B(N345));
XOR2X1 uut68 (.Y(N350),.A(N270),.B(N338));
XOR2X1 uut69 (.Y(N351),.A(N271),.B(N339));
XOR2X1 uut70 (.Y(N352),.A(N272),.B(N340));
XOR2X1 uut71 (.Y(N353),.A(N273),.B(N341));
XOR2X1 uut72 (.Y(N354),.A(N314),.B(N346));
XOR2X1 uut73 (.Y(N367),.A(N315),.B(N347));
XOR2X1 uut74 (.Y(N380),.A(N316),.B(N348));
XOR2X1 uut75 (.Y(N393),.A(N317),.B(N349));
XOR2X1 uut76 (.Y(N406),.A(N318),.B(N350));
XOR2X1 uut77 (.Y(N419),.A(N319),.B(N351));
XOR2X1 uut78 (.Y(N432),.A(N320),.B(N352));
XOR2X1 uut79 (.Y(N445),.A(N321),.B(N353));
INVX1 uut80 (.Y(N554),.A(N354fo0));
INVX1 uut81 (.Y(N555),.A(N367fo0));
INVX1 uut82 (.Y(N556),.A(N380fo0));
INVX1 uut83 (.Y(N557),.A(N354fo1));
INVX1 uut84 (.Y(N558),.A(N367fo1));
INVX1 uut85 (.Y(N559),.A(N393fo0));
INVX1 uut86 (.Y(N560),.A(N354fo2));
INVX1 uut87 (.Y(N561),.A(N380fo1));
INVX1 uut88 (.Y(N562),.A(N393fo1));
INVX1 uut89 (.Y(N563),.A(N367fo2));
INVX1 uut90 (.Y(N564),.A(N380fo2));
INVX1 uut91 (.Y(N565),.A(N393fo2));
INVX1 uut92 (.Y(N566),.A(N419fo0));
INVX1 uut93 (.Y(N567),.A(N445fo0));
INVX1 uut94 (.Y(N568),.A(N419fo1));
INVX1 uut95 (.Y(N569),.A(N432fo0));
INVX1 uut96 (.Y(N570),.A(N406fo0));
INVX1 uut97 (.Y(N571),.A(N445fo1));
INVX1 uut98 (.Y(N572),.A(N406fo1));
INVX1 uut99 (.Y(N573),.A(N432fo1));
INVX1 uut100 (.Y(N574),.A(N406fo2));
INVX1 uut101 (.Y(N575),.A(N419fo2));
INVX1 uut102 (.Y(N576),.A(N432fo2));
INVX1 uut103 (.Y(N577),.A(N406fo3));
INVX1 uut104 (.Y(N578),.A(N419fo3));
INVX1 uut105 (.Y(N579),.A(N445fo2));
INVX1 uut106 (.Y(N580),.A(N406fo4));
INVX1 uut107 (.Y(N581),.A(N432fo3));
INVX1 uut108 (.Y(N582),.A(N445fo3));
INVX1 uut109 (.Y(N583),.A(N419fo4));
INVX1 uut110 (.Y(N584),.A(N432fo4));
INVX1 uut111 (.Y(N585),.A(N445fo4));
INVX1 uut112 (.Y(N586),.A(N367fo3));
INVX1 uut113 (.Y(N587),.A(N393fo3));
INVX1 uut114 (.Y(N588),.A(N367fo4));
INVX1 uut115 (.Y(N589),.A(N380fo3));
INVX1 uut116 (.Y(N590),.A(N354fo3));
INVX1 uut117 (.Y(N591),.A(N393fo4));
INVX1 uut118 (.Y(N592),.A(N354fo4));
INVX1 uut119 (.Y(N593),.A(N380fo4));
AND2X1 uut120 (.Y(ttmp1),.A(N556),.B(N393fo5));
AND2X1 uut121 (.Y(ttmp2),.A(N554),.B(ttmp1));
AND2X1 uut122 (.Y(N594),.A(N555),.B(ttmp2));
AND2X1 uut123 (.Y(ttmp4),.A(N380fo5),.B(N559));
AND2X1 uut124 (.Y(ttmp5),.A(N557),.B(ttmp4));
AND2X1 uut125 (.Y(N595),.A(N558),.B(ttmp5));
AND2X1 uut126 (.Y(ttmp7),.A(N561),.B(N562));
AND2X1 uut127 (.Y(ttmp8),.A(N560),.B(ttmp7));
AND2X1 uut128 (.Y(N596),.A(N367fo5),.B(ttmp8));
AND2X1 uut129 (.Y(ttmp10),.A(N564),.B(N565));
AND2X1 uut130 (.Y(ttmp11),.A(N354fo5),.B(ttmp10));
AND2X1 uut131 (.Y(N597),.A(N563),.B(ttmp11));
AND2X1 uut132 (.Y(ttmp13),.A(N576),.B(N445fo5));
AND2X1 uut133 (.Y(ttmp14),.A(N574),.B(ttmp13));
AND2X1 uut134 (.Y(N598),.A(N575),.B(ttmp14));
AND2X1 uut135 (.Y(ttmp16),.A(N432fo5),.B(N579));
AND2X1 uut136 (.Y(ttmp17),.A(N577),.B(ttmp16));
AND2X1 uut137 (.Y(N599),.A(N578),.B(ttmp17));
AND2X1 uut138 (.Y(ttmp19),.A(N581),.B(N582));
AND2X1 uut139 (.Y(ttmp20),.A(N580),.B(ttmp19));
AND2X1 uut140 (.Y(N600),.A(N419fo5),.B(ttmp20));
AND2X1 uut141 (.Y(ttmp22),.A(N584),.B(N585));
AND2X1 uut142 (.Y(ttmp23),.A(N406fo5),.B(ttmp22));
AND2X1 uut143 (.Y(N601),.A(N583),.B(ttmp23));
OR2X1 uut144 (.Y(ttmp25),.A(N596),.B(N597));
OR2X1 uut145 (.Y(ttmp26),.A(N594),.B(ttmp25));
OR2X1 uut146 (.Y(N602),.A(N595),.B(ttmp26));
OR2X1 uut147 (.Y(ttmp28),.A(N600),.B(N601));
OR2X1 uut148 (.Y(ttmp29),.A(N598),.B(ttmp28));
OR2X1 uut149 (.Y(N607),.A(N599),.B(ttmp29));
AND2X1 uut150 (.Y(ttmp31),.A(N567),.B(N602fo0));
AND2X1 uut151 (.Y(ttmp32),.A(N406fo6),.B(ttmp31));
AND2X1 uut152 (.Y(ttmp33),.A(N566),.B(ttmp32));
AND2X1 uut153 (.Y(N620),.A(N432fo6),.B(ttmp33));
AND2X1 uut154 (.Y(ttmp35),.A(N445fo6),.B(N602fo1));
AND2X1 uut155 (.Y(ttmp36),.A(N406fo7),.B(ttmp35));
AND2X1 uut156 (.Y(ttmp37),.A(N568),.B(ttmp36));
AND2X1 uut157 (.Y(N625),.A(N569),.B(ttmp37));
AND2X1 uut158 (.Y(ttmp39),.A(N571),.B(N602fo2));
AND2X1 uut159 (.Y(ttmp40),.A(N570),.B(ttmp39));
AND2X1 uut160 (.Y(ttmp41),.A(N419fo6),.B(ttmp40));
AND2X1 uut161 (.Y(N630),.A(N432fo7),.B(ttmp41));
AND2X1 uut162 (.Y(ttmp43),.A(N445fo7),.B(N602fo3));
AND2X1 uut163 (.Y(ttmp44),.A(N572),.B(ttmp43));
AND2X1 uut164 (.Y(ttmp45),.A(N419fo7),.B(ttmp44));
AND2X1 uut165 (.Y(N635),.A(N573),.B(ttmp45));
AND2X1 uut166 (.Y(ttmp47),.A(N587),.B(N607fo0));
AND2X1 uut167 (.Y(ttmp48),.A(N354fo6),.B(ttmp47));
AND2X1 uut168 (.Y(ttmp49),.A(N586),.B(ttmp48));
AND2X1 uut169 (.Y(N640),.A(N380fo6),.B(ttmp49));
AND2X1 uut170 (.Y(ttmp51),.A(N393fo6),.B(N607fo1));
AND2X1 uut171 (.Y(ttmp52),.A(N354fo7),.B(ttmp51));
AND2X1 uut172 (.Y(ttmp53),.A(N588),.B(ttmp52));
AND2X1 uut173 (.Y(N645),.A(N589),.B(ttmp53));
AND2X1 uut174 (.Y(ttmp55),.A(N591),.B(N607fo2));
AND2X1 uut175 (.Y(ttmp56),.A(N590),.B(ttmp55));
AND2X1 uut176 (.Y(ttmp57),.A(N367fo6),.B(ttmp56));
AND2X1 uut177 (.Y(N650),.A(N380fo7),.B(ttmp57));
AND2X1 uut178 (.Y(ttmp59),.A(N393fo7),.B(N607fo3));
AND2X1 uut179 (.Y(ttmp60),.A(N592),.B(ttmp59));
AND2X1 uut180 (.Y(ttmp61),.A(N367fo7),.B(ttmp60));
AND2X1 uut181 (.Y(N655),.A(N593),.B(ttmp61));
AND2X1 uut182 (.Y(N692),.A(N354fo8),.B(N620fo0));
AND2X1 uut183 (.Y(N693),.A(N367fo8),.B(N620fo1));
AND2X1 uut184 (.Y(N694),.A(N380fo8),.B(N620fo2));
AND2X1 uut185 (.Y(N695),.A(N393fo8),.B(N620fo3));
AND2X1 uut186 (.Y(N696),.A(N354fo9),.B(N625fo0));
AND2X1 uut187 (.Y(N697),.A(N367fo9),.B(N625fo1));
AND2X1 uut188 (.Y(N698),.A(N380fo9),.B(N625fo2));
AND2X1 uut189 (.Y(N699),.A(N393fo9),.B(N625fo3));
AND2X1 uut190 (.Y(N700),.A(N354fo10),.B(N630fo0));
AND2X1 uut191 (.Y(N701),.A(N367fo10),.B(N630fo1));
AND2X1 uut192 (.Y(N702),.A(N380fo10),.B(N630fo2));
AND2X1 uut193 (.Y(N703),.A(N393fo10),.B(N630fo3));
AND2X1 uut194 (.Y(N704),.A(N354fo11),.B(N635fo0));
AND2X1 uut195 (.Y(N705),.A(N367fo11),.B(N635fo1));
AND2X1 uut196 (.Y(N706),.A(N380fo11),.B(N635fo2));
AND2X1 uut197 (.Y(N707),.A(N393fo11),.B(N635fo3));
AND2X1 uut198 (.Y(N708),.A(N406fo8),.B(N640fo0));
AND2X1 uut199 (.Y(N709),.A(N419fo8),.B(N640fo1));
AND2X1 uut200 (.Y(N710),.A(N432fo8),.B(N640fo2));
AND2X1 uut201 (.Y(N711),.A(N445fo8),.B(N640fo3));
AND2X1 uut202 (.Y(N712),.A(N406fo9),.B(N645fo0));
AND2X1 uut203 (.Y(N713),.A(N419fo9),.B(N645fo1));
AND2X1 uut204 (.Y(N714),.A(N432fo9),.B(N645fo2));
AND2X1 uut205 (.Y(N715),.A(N445fo9),.B(N645fo3));
AND2X1 uut206 (.Y(N716),.A(N406fo10),.B(N650fo0));
AND2X1 uut207 (.Y(N717),.A(N419fo10),.B(N650fo1));
AND2X1 uut208 (.Y(N718),.A(N432fo10),.B(N650fo2));
AND2X1 uut209 (.Y(N719),.A(N445fo10),.B(N650fo3));
AND2X1 uut210 (.Y(N720),.A(N406fo11),.B(N655fo0));
AND2X1 uut211 (.Y(N721),.A(N419fo11),.B(N655fo1));
AND2X1 uut212 (.Y(N722),.A(N432fo11),.B(N655fo2));
AND2X1 uut213 (.Y(N723),.A(N445fo11),.B(N655fo3));
XOR2X1 uut214 (.Y(N724),.A(N1fo2),.B(N692));
XOR2X1 uut215 (.Y(N725),.A(N5fo2),.B(N693));
XOR2X1 uut216 (.Y(N726),.A(N9fo2),.B(N694));
XOR2X1 uut217 (.Y(N727),.A(N13fo2),.B(N695));
XOR2X1 uut218 (.Y(N728),.A(N17fo2),.B(N696));
XOR2X1 uut219 (.Y(N729),.A(N21fo2),.B(N697));
XOR2X1 uut220 (.Y(N730),.A(N25fo2),.B(N698));
XOR2X1 uut221 (.Y(N731),.A(N29fo2),.B(N699));
XOR2X1 uut222 (.Y(N732),.A(N33fo2),.B(N700));
XOR2X1 uut223 (.Y(N733),.A(N37fo2),.B(N701));
XOR2X1 uut224 (.Y(N734),.A(N41fo2),.B(N702));
XOR2X1 uut225 (.Y(N735),.A(N45fo2),.B(N703));
XOR2X1 uut226 (.Y(N736),.A(N49fo2),.B(N704));
XOR2X1 uut227 (.Y(N737),.A(N53fo2),.B(N705));
XOR2X1 uut228 (.Y(N738),.A(N57fo2),.B(N706));
XOR2X1 uut229 (.Y(N739),.A(N61fo2),.B(N707));
XOR2X1 uut230 (.Y(N740),.A(N65fo2),.B(N708));
XOR2X1 uut231 (.Y(N741),.A(N69fo2),.B(N709));
XOR2X1 uut232 (.Y(N742),.A(N73fo2),.B(N710));
XOR2X1 uut233 (.Y(N743),.A(N77fo2),.B(N711));
XOR2X1 uut234 (.Y(N744),.A(N81fo2),.B(N712));
XOR2X1 uut235 (.Y(N745),.A(N85fo2),.B(N713));
XOR2X1 uut236 (.Y(N746),.A(N89fo2),.B(N714));
XOR2X1 uut237 (.Y(N747),.A(N93fo2),.B(N715));
XOR2X1 uut238 (.Y(N748),.A(N97fo2),.B(N716));
XOR2X1 uut239 (.Y(N749),.A(N101fo2),.B(N717));
XOR2X1 uut240 (.Y(N750),.A(N105fo2),.B(N718));
XOR2X1 uut241 (.Y(N751),.A(N109fo2),.B(N719));
XOR2X1 uut242 (.Y(N752),.A(N113fo2),.B(N720));
XOR2X1 uut243 (.Y(N753),.A(N117fo2),.B(N721));
XOR2X1 uut244 (.Y(N754),.A(N121fo2),.B(N722));
XOR2X1 uut245 (.Y(N755),.A(N125fo2),.B(N723));
fanout3 uut_fo0 (.A(N1),.Y1(N1fo0),.Y2(N1fo1),.Y3(N1fo2));
fanout3 uut_fo1 (.A(N5),.Y1(N5fo0),.Y2(N5fo1),.Y3(N5fo2));
fanout3 uut_fo2 (.A(N9),.Y1(N9fo0),.Y2(N9fo1),.Y3(N9fo2));
fanout3 uut_fo3 (.A(N13),.Y1(N13fo0),.Y2(N13fo1),.Y3(N13fo2));
fanout3 uut_fo4 (.A(N17),.Y1(N17fo0),.Y2(N17fo1),.Y3(N17fo2));
fanout3 uut_fo5 (.A(N21),.Y1(N21fo0),.Y2(N21fo1),.Y3(N21fo2));
fanout3 uut_fo6 (.A(N25),.Y1(N25fo0),.Y2(N25fo1),.Y3(N25fo2));
fanout3 uut_fo7 (.A(N29),.Y1(N29fo0),.Y2(N29fo1),.Y3(N29fo2));
fanout3 uut_fo8 (.A(N33),.Y1(N33fo0),.Y2(N33fo1),.Y3(N33fo2));
fanout3 uut_fo9 (.A(N37),.Y1(N37fo0),.Y2(N37fo1),.Y3(N37fo2));
fanout3 uut_fo10 (.A(N41),.Y1(N41fo0),.Y2(N41fo1),.Y3(N41fo2));
fanout3 uut_fo11 (.A(N45),.Y1(N45fo0),.Y2(N45fo1),.Y3(N45fo2));
fanout3 uut_fo12 (.A(N49),.Y1(N49fo0),.Y2(N49fo1),.Y3(N49fo2));
fanout3 uut_fo13 (.A(N53),.Y1(N53fo0),.Y2(N53fo1),.Y3(N53fo2));
fanout3 uut_fo14 (.A(N57),.Y1(N57fo0),.Y2(N57fo1),.Y3(N57fo2));
fanout3 uut_fo15 (.A(N61),.Y1(N61fo0),.Y2(N61fo1),.Y3(N61fo2));
fanout3 uut_fo16 (.A(N65),.Y1(N65fo0),.Y2(N65fo1),.Y3(N65fo2));
fanout3 uut_fo17 (.A(N69),.Y1(N69fo0),.Y2(N69fo1),.Y3(N69fo2));
fanout3 uut_fo18 (.A(N73),.Y1(N73fo0),.Y2(N73fo1),.Y3(N73fo2));
fanout3 uut_fo19 (.A(N77),.Y1(N77fo0),.Y2(N77fo1),.Y3(N77fo2));
fanout3 uut_fo20 (.A(N81),.Y1(N81fo0),.Y2(N81fo1),.Y3(N81fo2));
fanout3 uut_fo21 (.A(N85),.Y1(N85fo0),.Y2(N85fo1),.Y3(N85fo2));
fanout3 uut_fo22 (.A(N89),.Y1(N89fo0),.Y2(N89fo1),.Y3(N89fo2));
fanout3 uut_fo23 (.A(N93),.Y1(N93fo0),.Y2(N93fo1),.Y3(N93fo2));
fanout3 uut_fo24 (.A(N97),.Y1(N97fo0),.Y2(N97fo1),.Y3(N97fo2));
fanout3 uut_fo25 (.A(N101),.Y1(N101fo0),.Y2(N101fo1),.Y3(N101fo2));
fanout3 uut_fo26 (.A(N105),.Y1(N105fo0),.Y2(N105fo1),.Y3(N105fo2));
fanout3 uut_fo27 (.A(N109),.Y1(N109fo0),.Y2(N109fo1),.Y3(N109fo2));
fanout3 uut_fo28 (.A(N113),.Y1(N113fo0),.Y2(N113fo1),.Y3(N113fo2));
fanout3 uut_fo29 (.A(N117),.Y1(N117fo0),.Y2(N117fo1),.Y3(N117fo2));
fanout3 uut_fo30 (.A(N121),.Y1(N121fo0),.Y2(N121fo1),.Y3(N121fo2));
fanout3 uut_fo31 (.A(N125),.Y1(N125fo0),.Y2(N125fo1),.Y3(N125fo2));
fanout8 uut_fo40 (.A(N137),.Y1(N137fo0),.Y2(N137fo1),.Y3(N137fo2),.Y4(N137fo3),.Y5(N137fo4),.Y6(N137fo5),.Y7(N137fo6),.Y8(N137fo7));
fanout12 uut_fo_w4 (.A(N445),.Y1(N445fo0),.Y2(N445fo1),.Y3(N445fo2),.Y4(N445fo3),.Y5(N445fo4),.Y6(N445fo5),.Y7(N445fo6),.Y8(N445fo7),.Y9(N445fo8),.Y10(N445fo9),.Y11(N445fo10),.Y12(N445fo11));
fanout4 uut_fo_w5 (.A(N630),.Y1(N630fo0),.Y2(N630fo1),.Y3(N630fo2),.Y4(N630fo3));
fanout4 uut_fo_w28 (.A(N602),.Y1(N602fo0),.Y2(N602fo1),.Y3(N602fo2),.Y4(N602fo3));
fanout4 uut_fo_w40 (.A(N607),.Y1(N607fo0),.Y2(N607fo1),.Y3(N607fo2),.Y4(N607fo3));
fanout4 uut_fo_w49 (.A(N625),.Y1(N625fo0),.Y2(N625fo1),.Y3(N625fo2),.Y4(N625fo3));
fanout2 uut_fo_w68 (.A(N308),.Y1(N308fo0),.Y2(N308fo1));
fanout2 uut_fo_w73 (.A(N293),.Y1(N293fo0),.Y2(N293fo1));
fanout12 uut_fo_w77 (.A(N406),.Y1(N406fo0),.Y2(N406fo1),.Y3(N406fo2),.Y4(N406fo3),.Y5(N406fo4),.Y6(N406fo5),.Y7(N406fo6),.Y8(N406fo7),.Y9(N406fo8),.Y10(N406fo9),.Y11(N406fo10),.Y12(N406fo11));
fanout2 uut_fo_w105 (.A(N302),.Y1(N302fo0),.Y2(N302fo1));
fanout2 uut_fo_w116 (.A(N299),.Y1(N299fo0),.Y2(N299fo1));
fanout12 uut_fo_w124 (.A(N432),.Y1(N432fo0),.Y2(N432fo1),.Y3(N432fo2),.Y4(N432fo3),.Y5(N432fo4),.Y6(N432fo5),.Y7(N432fo6),.Y8(N432fo7),.Y9(N432fo8),.Y10(N432fo9),.Y11(N432fo10),.Y12(N432fo11));
fanout4 uut_fo_w127 (.A(N635),.Y1(N635fo0),.Y2(N635fo1),.Y3(N635fo2),.Y4(N635fo3));
fanout4 uut_fo_w134 (.A(N645),.Y1(N645fo0),.Y2(N645fo1),.Y3(N645fo2),.Y4(N645fo3));
fanout2 uut_fo_w135 (.A(N296),.Y1(N296fo0),.Y2(N296fo1));
fanout4 uut_fo_w152 (.A(N655),.Y1(N655fo0),.Y2(N655fo1),.Y3(N655fo2),.Y4(N655fo3));
fanout4 uut_fo_w154 (.A(N620),.Y1(N620fo0),.Y2(N620fo1),.Y3(N620fo2),.Y4(N620fo3));
fanout12 uut_fo_w155 (.A(N393),.Y1(N393fo0),.Y2(N393fo1),.Y3(N393fo2),.Y4(N393fo3),.Y5(N393fo4),.Y6(N393fo5),.Y7(N393fo6),.Y8(N393fo7),.Y9(N393fo8),.Y10(N393fo9),.Y11(N393fo10),.Y12(N393fo11));
fanout4 uut_fo_w156 (.A(N650),.Y1(N650fo0),.Y2(N650fo1),.Y3(N650fo2),.Y4(N650fo3));
fanout12 uut_fo_w157 (.A(N367),.Y1(N367fo0),.Y2(N367fo1),.Y3(N367fo2),.Y4(N367fo3),.Y5(N367fo4),.Y6(N367fo5),.Y7(N367fo6),.Y8(N367fo7),.Y9(N367fo8),.Y10(N367fo9),.Y11(N367fo10),.Y12(N367fo11));
fanout2 uut_fo_w167 (.A(N311),.Y1(N311fo0),.Y2(N311fo1));
fanout2 uut_fo_w183 (.A(N305),.Y1(N305fo0),.Y2(N305fo1));
fanout12 uut_fo_w188 (.A(N419),.Y1(N419fo0),.Y2(N419fo1),.Y3(N419fo2),.Y4(N419fo3),.Y5(N419fo4),.Y6(N419fo5),.Y7(N419fo6),.Y8(N419fo7),.Y9(N419fo8),.Y10(N419fo9),.Y11(N419fo10),.Y12(N419fo11));
fanout12 uut_fo_w192 (.A(N354),.Y1(N354fo0),.Y2(N354fo1),.Y3(N354fo2),.Y4(N354fo3),.Y5(N354fo4),.Y6(N354fo5),.Y7(N354fo6),.Y8(N354fo7),.Y9(N354fo8),.Y10(N354fo9),.Y11(N354fo10),.Y12(N354fo11));
fanout12 uut_fo_w196 (.A(N380),.Y1(N380fo0),.Y2(N380fo1),.Y3(N380fo2),.Y4(N380fo3),.Y5(N380fo4),.Y6(N380fo5),.Y7(N380fo6),.Y8(N380fo7),.Y9(N380fo8),.Y10(N380fo9),.Y11(N380fo10),.Y12(N380fo11));
fanout4 uut_fo_w203 (.A(N640),.Y1(N640fo0),.Y2(N640fo1),.Y3(N640fo2),.Y4(N640fo3));
fanout2 uut_fo_w208 (.A(N290),.Y1(N290fo0),.Y2(N290fo1));
endmodule